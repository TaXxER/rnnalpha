20000 4
7 3 0 3 1 3 1 3
2 3 3
5 3 2 0 3 0
4 3 0 1 0
7 3 3 0 0 1 3 0
2 3 1
4 3 0 3 3
5 3 0 3 1 3
23 3 1 3 0 2 0 3 1 2 0 3 0 2 0 1 0 3 0 1 0 3 3 3
2 3 0
2 3 3
17 3 3 0 1 1 1 1 1 1 1 1 2 0 3 0 2 1
3 3 1 3
27 3 0 1 2 0 3 1 2 2 1 3 0 0 3 3 1 0 1 3 3 1 3 0 3 0 2 3
4 3 1 2 0
2 3 3
3 3 3 3
3 3 0 1
22 3 3 1 3 3 1 3 3 3 1 3 3 3 0 0 3 0 0 0 3 3 1
3 3 0 3
17 3 0 3 1 0 1 3 3 2 0 1 3 1 3 2 0 3
35 3 3 0 2 3 1 3 0 3 0 3 1 1 3 3 0 3 0 1 0 1 3 3 1 2 2 0 3 0 1 1 1 1 3 3
3 3 0 3
16 3 0 3 3 3 0 2 3 0 2 0 3 1 3 1 2
11 3 0 3 1 3 0 3 0 1 3 3
4 3 1 0 3
3 3 3 1
5 3 3 1 3 3
3 3 0 2
15 3 0 2 1 1 3 1 1 3 3 0 3 0 1 2
13 3 0 3 1 2 2 3 2 0 2 0 3 0
2 3 3
3 3 3 0
18 3 1 1 3 0 2 1 2 2 2 0 0 3 0 1 0 0 3
13 3 1 3 2 0 0 0 1 1 1 2 3 0
3 3 0 3
3 3 3 0
5 3 3 1 0 0
8 3 3 2 0 0 1 3 0
3 3 0 2
4 3 1 3 0
3 3 0 3
16 3 3 0 1 1 1 1 1 1 1 0 3 0 1 2 3
2 3 3
3 3 1 2
7 3 3 1 3 3 1 3
4 3 0 2 3
2 3 0
5 3 0 1 3 1
7 3 0 3 1 2 1 3
8 3 1 1 1 1 1 1 1
3 3 1 3
31 3 0 3 0 0 2 0 2 0 3 0 1 3 3 1 2 1 2 0 3 1 0 1 3 3 1 1 3 3 2 0
24 3 0 0 0 2 3 1 2 3 1 0 2 3 1 3 0 0 1 3 3 0 0 0 2
19 3 0 3 3 1 3 3 0 3 0 1 2 3 0 3 0 3 0 2
17 3 0 1 3 3 0 3 0 1 3 3 3 1 3 3 3 0
19 3 3 0 1 2 0 3 0 1 1 3 0 3 0 3 0 1 3 1
3 3 1 3
11 3 0 3 0 0 3 1 2 2 1 3
7 3 0 3 1 3 0 3
19 3 1 3 0 2 0 2 3 0 2 1 1 1 3 0 2 0 3 0
11 3 1 3 0 0 0 1 0 2 3 2
3 3 0 3
10 3 0 3 1 2 1 3 2 0 3
14 3 0 3 1 2 2 0 3 0 1 3 3 0 2
2 3 3
8 3 3 1 3 3 1 3 0
17 3 0 3 0 0 3 1 0 1 3 3 0 2 0 1 3 0
1 3
24 3 0 3 0 0 3 0 1 3 3 3 0 1 2 0 2 2 1 1 0 2 1 0 3
5 3 3 1 3 3
26 3 0 3 1 2 1 1 1 1 1 3 0 2 3 0 0 1 3 0 0 1 3 1 1 3 2
4 3 2 0 3
3 3 1 3
4 3 1 3 0
2 3 3
3 3 1 2
6 3 3 0 2 3 3
8 3 1 1 3 2 0 3 3
8 3 0 3 0 1 3 3 2
13 3 2 2 0 1 2 2 3 1 1 3 0 2
3 3 0 3
24 3 3 1 3 3 0 3 0 3 3 3 0 1 1 3 1 0 1 2 1 3 3 0 3
4 3 0 2 3
2 3 3
2 3 3
4 3 1 2 0
4 3 1 1 1
3 3 0 3
26 3 3 0 2 0 3 0 2 0 3 3 1 3 3 0 2 3 0 1 3 2 0 1 3 1 1
6 3 3 1 0 1 3
4 3 2 2 0
12 3 0 3 0 3 0 1 3 3 0 1 2
14 3 0 2 0 0 0 1 3 0 2 0 3 0 2
6 3 0 3 1 0 2
7 3 1 2 1 3 3 3
3 3 1 2
3 3 3 0
5 3 0 1 1 3
3 3 0 3
5 3 0 3 0 1
4 3 0 2 3
1 3
19 3 0 2 3 0 0 0 3 3 3 0 1 3 3 3 0 0 0 1
1 3
1 3
4 3 3 1 1
5 3 0 3 1 3
3 3 0 3
5 3 1 2 1 1
18 3 3 0 2 0 3 1 2 1 1 1 2 3 2 3 1 2 1
3 3 1 3
3 3 3 0
3 3 3 0
3 3 1 2
4 3 0 2 3
3 3 1 3
4 3 0 2 0
2 3 0
12 3 0 3 3 1 0 3 1 2 1 1 1
7 3 0 3 0 0 3 0
5 3 0 1 3 3
3 3 0 3
2 3 3
5 3 0 2 3 0
7 3 0 3 1 1 3 3
3 3 1 3
6 3 0 3 0 0 3
2 3 3
16 3 3 1 3 1 3 0 1 2 0 3 0 1 3 3 3
12 3 3 0 1 1 1 1 1 1 2 0 3
4 3 1 1 3
5 3 3 1 3 3
6 3 1 0 3 1 2
8 3 0 3 1 3 3 0 2
1 3
3 3 1 3
3 3 1 3
7 3 1 3 0 0 3 0
18 3 1 2 0 1 3 3 0 2 3 1 3 0 0 0 0 0 1
2 3 0
7 3 0 3 0 2 0 3
5 3 0 1 2 3
5 3 3 2 0 2
21 3 0 3 0 1 3 3 1 3 0 2 3 1 1 0 0 1 2 1 1 3
3 3 0 1
1 3
3 3 0 3
1 3
3 3 1 1
27 3 0 3 1 0 2 0 0 2 1 1 2 2 0 2 3 1 3 3 3 1 3 3 0 3 0 3
3 3 0 3
7 3 0 3 1 2 0 3
22 3 0 3 1 2 2 3 1 3 1 3 0 1 1 2 0 1 0 0 1 0 2
7 3 3 0 2 3 3 0
5 3 0 3 0 2
4 3 0 3 0
4 3 1 1 3
3 3 0 3
2 3 3
4 3 3 3 0
5 3 1 3 2 1
3 3 3 0
3 3 0 3
2 3 3
1 3
3 3 1 3
6 3 0 3 0 2 0
2 3 3
2 3 3
2 3 2
8 3 0 3 0 1 1 3 3
3 3 0 3
2 3 3
14 3 0 2 3 1 3 3 0 1 3 3 1 3 3
9 3 0 3 1 2 1 0 0 3
2 3 3
7 3 0 1 3 3 3 0
3 3 1 3
6 3 1 3 1 3 1
6 3 1 3 0 2 1
3 3 1 3
4 3 1 1 3
5 3 0 1 0 0
6 3 3 0 0 3 1
2 3 3
4 3 1 2 0
4 3 0 2 3
10 3 0 3 0 1 3 3 0 2 3
8 3 0 3 0 3 0 1 3
4 3 1 3 0
4 3 2 0 3
1 3
2 3 3
5 3 0 3 3 0
3 3 0 3
4 3 3 2 3
3 3 3 2
1 3
13 3 0 3 0 3 0 1 3 3 0 3 0 3
3 3 0 3
4 3 1 1 3
7 3 0 3 1 3 1 3
4 3 1 1 3
4 3 0 2 3
3 3 3 0
3 3 1 3
9 3 1 1 3 1 1 1 1 1
4 3 0 2 3
4 3 0 3 0
4 3 3 0 2
9 3 3 1 3 3 0 1 0 3
5 3 3 0 2 2
6 3 0 3 1 0 2
13 3 3 3 0 0 1 3 0 1 2 1 3 0
19 3 0 3 1 3 1 1 3 0 1 3 1 3 3 3 0 2 0 3
10 3 0 3 0 1 3 3 1 2 2
4 3 3 1 0
10 3 2 0 1 3 0 0 1 3 0
12 3 1 1 3 0 1 1 0 1 3 2 3
2 3 3
2 3 3
4 3 3 1 3
3 3 3 0
1 3
1 3
2 3 3
13 3 0 3 1 2 2 0 3 0 3 1 0 2
5 3 0 2 3 0
5 3 0 3 1 3
10 3 1 3 1 2 0 2 3 3 0
9 3 0 3 0 1 0 1 3 0
3 3 0 3
4 3 0 2 3
2 3 0
4 3 0 2 3
8 3 0 3 0 0 1 0 0
5 3 0 3 1 2
2 3 3
14 3 0 2 2 1 2 0 2 3 1 1 1 1 1
5 3 0 3 0 0
9 3 0 3 0 2 3 3 3 0
6 3 3 0 1 2 3
4 3 1 1 2
3 3 3 0
4 3 0 3 3
11 3 3 1 3 3 3 1 2 3 0 0
14 3 0 2 3 0 1 0 0 0 3 1 2 3 0
12 3 1 2 0 2 3 1 1 1 3 1 3
3 3 0 3
7 3 3 1 3 3 0 3
9 3 3 1 3 3 3 1 3 1
1 3
11 3 0 3 3 1 3 3 3 2 3 0
4 3 3 0 3
11 3 3 1 3 3 0 3 0 0 3 0
4 3 0 2 3
7 3 0 3 0 1 3 3
10 3 3 1 1 3 0 1 2 1 0
3 3 3 0
12 3 3 0 2 0 3 0 1 2 0 2 3
8 3 3 0 1 0 1 2 3
11 3 0 3 0 3 1 2 0 2 1 0
7 3 0 1 2 3 3 0
7 3 0 3 1 2 3 0
6 3 1 3 0 0 0
4 3 3 0 0
14 3 3 0 2 1 1 1 1 1 1 1 3 0 0
3 3 0 3
14 3 0 0 2 3 3 2 1 0 1 3 3 0 3
5 3 0 1 2 3
15 3 1 1 3 3 3 1 3 0 1 2 3 0 2 1
7 3 1 2 1 1 1 3
4 3 0 3 3
30 3 1 1 1 1 3 3 2 1 3 2 1 2 3 1 3 3 1 3 0 0 0 3 2 3 3 0 1 2 3
13 3 1 0 3 3 3 1 3 3 0 1 3 3
6 3 1 3 0 1 1
3 3 0 3
13 3 0 3 0 1 3 3 1 3 0 2 0 2
6 3 3 0 2 0 3
19 3 3 0 2 2 0 3 1 3 3 1 3 0 2 0 1 3 3 0
31 3 0 3 1 2 3 0 0 1 3 1 3 0 1 1 2 2 0 3 0 1 3 3 0 1 1 0 1 3 0 3
17 3 1 1 1 3 0 2 3 0 3 1 2 0 1 3 3 3
2 3 3
3 3 0 3
3 3 3 0
14 3 1 3 0 2 1 0 3 3 0 1 1 1 1
4 3 0 3 0
8 3 0 3 0 2 0 1 3
15 3 3 1 3 3 1 2 1 3 2 1 2 3 0 0
18 3 3 0 0 1 3 0 2 2 0 3 1 1 1 1 2 2 3
3 3 3 0
7 3 0 3 1 2 1 1
10 3 0 2 3 0 3 1 2 3 0
3 3 1 3
12 3 0 3 1 2 1 1 1 1 1 0 1
1 3
6 3 3 0 1 1 0
10 3 0 3 1 2 1 3 3 3 3
6 3 1 1 1 1 3
3 3 0 3
2 3 3
4 3 3 0 1
2 3 3
31 3 1 1 3 1 0 3 3 1 3 1 0 0 1 1 3 0 1 3 2 2 1 0 1 3 3 3 2 1 0 3
6 3 0 3 1 2 3
5 3 0 1 3 3
8 3 0 3 0 2 0 0 0
3 3 3 0
5 3 0 3 0 2
8 3 3 1 3 3 0 3 0
14 3 0 2 3 0 1 3 0 2 0 3 1 2 3
15 3 0 3 3 3 0 1 2 0 3 0 1 1 1 3
9 3 0 3 0 1 3 3 0 3
9 3 3 1 3 3 1 3 3 3
10 3 0 3 0 1 0 0 2 0 3
10 3 3 1 2 1 3 2 1 2 1
3 3 0 3
3 3 0 3
9 3 0 3 1 2 0 3 0 2
4 3 0 2 3
3 3 3 0
4 3 0 3 0
4 3 3 2 0
5 3 0 3 0 3
8 3 1 0 3 3 0 2 3
6 3 0 3 3 1 3
14 3 1 1 3 0 0 0 0 3 2 1 1 1 0
25 3 0 3 1 0 2 1 2 0 0 0 1 1 3 2 1 1 2 3 0 3 2 0 1 3
2 3 0
3 3 0 3
11 3 3 1 3 3 3 0 2 2 0 3
3 3 1 3
9 3 1 3 0 1 0 1 3 0
5 3 3 1 3 3
5 3 0 3 0 2
2 3 3
11 3 0 3 3 1 0 1 3 3 0 3
3 3 1 3
9 3 0 3 0 1 2 1 1 3
21 3 3 1 3 1 3 0 1 2 3 0 3 3 0 3 0 1 1 3 1 3
6 3 0 3 1 1 3
3 3 1 3
7 3 0 3 0 3 3 0
10 3 3 3 3 3 0 3 3 0 3
24 3 0 3 1 3 3 1 3 3 0 2 0 0 3 1 3 0 2 1 3 0 0 0 1
9 3 1 3 0 2 2 0 1 3
15 3 3 1 1 3 2 0 3 0 1 1 1 1 1 1
4 3 3 0 1
3 3 0 2
2 3 3
10 3 3 0 3 3 0 1 3 3 3
9 3 1 2 0 1 2 0 3 3
12 3 3 0 0 0 1 1 2 3 0 0 0
8 3 0 3 0 1 3 3 0
7 3 2 0 3 0 0 0
6 3 0 3 0 0 3
3 3 1 1
6 3 1 1 1 1 3
7 3 3 0 1 1 3 1
6 3 0 3 0 1 2
14 3 0 3 0 3 1 3 3 1 3 3 3 3 0
10 3 0 3 3 1 3 1 3 0 0
25 3 3 1 1 1 1 1 3 1 3 0 0 0 1 0 3 3 0 1 0 1 3 3 0 1
3 3 3 0
3 3 3 0
6 3 0 3 0 1 2
11 3 3 1 2 0 1 2 0 3 1 3
12 3 1 0 1 0 1 3 3 3 2 3 2
7 3 3 0 0 1 3 0
5 3 0 2 3 1
3 3 0 3
6 3 3 0 2 1 2
3 3 3 1
4 3 1 1 1
5 3 0 3 1 2
7 3 0 2 0 0 2 2
2 3 3
9 3 3 0 0 3 3 3 0 0
4 3 0 3 0
10 3 1 2 0 2 1 3 0 0 0
6 3 0 2 3 0 3
8 3 0 3 3 1 0 3 3
2 3 3
15 3 0 3 0 3 0 1 3 3 0 3 0 1 2 1
10 3 0 3 1 1 3 0 0 3 3
3 3 0 3
13 3 3 0 0 3 0 0 1 2 0 3 0 2
2 3 3
6 3 0 1 3 3 3
2 3 3
2 3 3
9 3 0 2 3 0 2 0 3 3
4 3 3 0 1
3 3 3 0
10 3 0 3 0 3 1 2 0 0 2
7 3 0 3 1 3 2 3
4 3 0 2 3
2 3 3
3 3 2 3
26 3 0 3 0 1 2 3 3 1 3 3 1 2 1 2 3 1 3 3 0 3 1 3 1 3 3
12 3 3 0 3 3 3 3 1 2 3 1 0
7 3 3 0 2 1 3 0
2 3 3
7 3 3 1 3 3 1 2
7 3 0 3 0 1 0 3
7 3 3 1 1 1 1 1
12 3 0 3 0 1 3 1 1 0 1 3 3
3 3 0 3
37 3 0 3 0 1 2 1 1 3 3 3 3 3 3 0 1 3 1 2 0 2 0 0 1 3 3 0 3 0 0 3 1 0 1 2 3 0
6 3 0 3 0 0 3
9 3 1 2 0 0 0 3 0 0
7 3 0 3 0 1 2 0
1 3
2 3 3
15 3 3 2 1 0 1 2 1 1 1 1 3 0 0 3
3 3 3 3
2 3 3
6 3 1 0 3 3 3
2 3 3
9 3 1 3 0 2 0 1 3 3
5 3 1 1 2 3
6 3 0 2 3 0 0
7 3 0 3 1 2 1 1
10 3 1 1 1 1 1 3 3 3 0
6 3 0 3 0 2 3
8 3 1 0 0 0 1 0 3
6 3 0 3 0 1 0
2 3 3
10 3 3 1 3 3 0 1 2 1 3
2 3 3
5 3 1 3 0 0
5 3 0 3 0 2
12 3 1 1 3 1 3 0 1 1 1 1 3
3 3 3 0
8 3 3 0 1 1 2 0 1
4 3 1 3 0
5 3 1 1 3 3
5 3 0 3 0 3
5 3 0 2 1 3
9 3 0 3 1 2 0 3 1 1
4 3 0 3 0
18 3 3 2 0 1 3 3 3 0 1 0 3 3 0 3 1 3 3
6 3 3 3 1 3 0
5 3 3 1 1 1
3 3 0 3
2 3 0
9 3 1 3 0 2 0 3 0 3
8 3 0 2 2 0 3 0 2
2 3 3
4 3 1 1 3
5 3 0 3 0 3
7 3 0 3 0 2 0 0
5 3 0 3 1 3
3 3 0 3
8 3 0 3 0 3 0 2 0
3 3 0 3
2 3 3
9 3 0 3 3 0 2 1 2 3
6 3 0 2 3 0 2
8 3 0 3 0 3 1 2 3
6 3 0 3 0 3 0
12 3 1 3 0 1 1 1 2 0 2 1 3
5 3 3 1 3 3
6 3 1 1 1 1 3
13 3 1 3 1 3 3 3 1 3 3 0 3 3
11 3 0 3 0 1 3 3 3 3 0 1
9 3 0 3 3 0 0 1 3 0
9 3 3 3 2 0 2 1 2 3
7 3 3 3 3 1 3 3
8 3 2 0 1 3 0 1 0
21 3 0 3 1 0 0 3 1 3 1 1 3 0 1 3 0 2 2 2 3 0
31 3 0 3 1 0 1 3 3 0 3 0 1 3 3 0 1 3 3 1 1 1 1 1 1 1 1 1 1 3 1 3
1 3
22 3 3 0 1 1 1 1 2 0 3 3 2 3 1 3 3 0 3 3 1 3 3
2 3 1
15 3 0 0 3 2 2 3 1 3 3 1 3 0 0 0
12 3 0 3 0 3 0 0 3 0 1 3 3
13 3 0 3 3 1 3 3 0 1 2 1 1 3
3 3 0 3
1 3
10 3 0 3 1 0 1 3 3 1 3
1 3
4 3 0 3 0
5 3 0 3 0 3
3 3 1 0
5 3 0 3 0 3
3 3 3 0
10 3 3 0 1 2 0 3 1 2 3
4 3 0 0 2
2 3 2
3 3 0 3
11 3 3 1 3 3 1 3 0 2 0 3
8 3 0 3 0 3 0 1 2
7 3 2 3 0 1 3 3
7 3 3 0 1 1 1 1
2 3 3
17 3 3 3 1 3 2 2 0 3 1 3 0 3 1 0 1 3
1 3
14 3 0 3 3 1 3 3 0 1 3 3 3 0 0
10 3 0 3 1 3 0 3 0 1 0
14 3 1 1 3 0 2 0 2 3 3 1 1 3 0
8 3 0 1 2 1 1 2 0
7 3 3 1 1 0 3 3
3 3 0 1
10 3 1 3 0 0 0 1 0 2 0
4 3 0 2 3
6 3 3 1 3 3 0
2 3 3
8 3 0 3 1 0 1 3 3
8 3 0 3 0 1 2 0 3
5 3 0 3 0 2
1 3
2 3 3
8 3 3 0 0 0 1 2 1
17 3 3 1 2 3 3 0 1 2 3 0 1 1 3 2 0 3
13 3 0 3 0 1 2 3 1 3 1 3 0 0
6 3 0 3 0 0 1
10 3 1 3 1 3 0 0 2 3 0
2 3 3
13 3 0 3 3 1 0 0 1 3 0 0 1 1
4 3 0 3 1
2 3 3
5 3 1 1 1 1
15 3 3 1 0 0 1 3 3 3 0 2 0 1 2 1
2 3 1
16 3 0 2 3 0 1 2 0 3 1 0 1 0 1 0 0
2 3 3
23 3 3 0 2 0 3 0 1 3 3 2 3 0 0 3 3 0 3 1 3 3 3 2
3 3 1 3
13 3 3 2 1 1 2 1 1 1 1 3 2 3
10 3 3 2 3 1 1 1 1 1 3
5 3 0 3 3 3
7 3 1 3 0 2 0 2
11 3 3 0 1 1 2 3 1 3 3 1
4 3 0 3 0
9 3 0 3 0 1 1 1 1 1
8 3 0 2 3 1 3 3 3
5 3 3 1 3 3
29 3 3 1 3 3 1 2 1 2 0 3 0 2 0 3 0 1 3 2 1 2 1 3 0 2 0 1 0 0
5 3 0 2 3 1
7 3 3 0 2 0 2 3
9 3 3 1 1 3 2 2 1 3
2 3 3
2 3 3
10 3 3 0 0 1 3 0 0 1 3
7 3 1 3 3 0 0 0
12 3 2 0 3 0 1 1 0 1 2 1 3
13 3 0 3 1 0 1 2 2 3 3 1 2 2
3 3 1 3
5 3 1 3 1 3
2 3 3
4 3 3 0 2
2 3 3
3 3 3 0
1 3
10 3 1 1 3 0 0 3 3 3 3
4 3 0 1 0
2 3 3
2 3 3
3 3 0 3
6 3 0 3 3 3 3
6 3 1 1 3 3 3
8 3 3 0 0 0 0 1 3
4 3 2 0 3
17 3 2 0 0 3 0 1 1 3 2 1 3 1 1 1 1 3
12 3 3 3 2 0 2 0 3 0 0 1 2
2 3 3
8 3 0 1 2 1 0 1 3
27 3 2 2 0 0 1 3 1 1 1 1 1 1 1 1 3 0 1 3 3 3 3 1 3 3 3 0
5 3 0 3 3 0
9 3 0 3 1 3 1 1 2 0
20 3 0 3 1 2 2 3 0 1 1 2 3 0 1 2 3 2 2 2 3
4 3 3 0 1
9 3 2 2 0 1 2 0 2 3
3 3 3 2
2 3 3
1 3
5 3 3 1 0 0
5 3 1 1 3 0
3 3 3 0
2 3 3
10 3 1 0 3 2 0 2 0 3 1
3 3 1 3
4 3 0 2 0
6 3 3 3 0 0 0
4 3 3 0 0
8 3 1 1 3 3 3 0 3
4 3 3 0 1
2 3 3
7 3 0 3 0 1 0 0
11 3 3 1 3 3 3 1 3 3 3 0
6 3 3 0 2 0 3
2 3 3
2 3 0
8 3 0 3 0 3 1 3 3
3 3 3 0
11 3 3 1 3 2 3 3 3 3 0 1
3 3 0 3
6 3 3 2 0 0 2
10 3 3 0 2 0 3 1 3 0 3
2 3 3
18 3 0 3 0 2 1 3 1 3 1 1 2 3 0 1 1 2 3
8 3 0 3 0 2 1 1 3
5 3 1 1 1 3
6 3 0 3 3 1 3
3 3 0 3
4 3 3 2 3
20 3 0 3 0 1 2 0 1 2 1 3 0 1 2 0 3 0 2 1 0
2 3 3
2 3 3
4 3 0 3 0
12 3 0 3 0 0 1 2 3 1 3 3 3
4 3 1 0 0
1 3
10 3 0 2 3 1 0 2 3 3 3
14 3 3 0 1 1 1 2 0 3 1 3 3 0 0
3 3 3 0
23 3 3 1 2 3 0 3 0 3 0 1 3 3 0 1 2 1 2 0 3 0 2 0
4 3 3 3 0
2 3 3
3 3 1 3
11 3 1 3 0 2 1 1 3 1 3 0
9 3 0 3 1 0 1 3 3 3
6 3 1 0 1 3 0
2 3 3
1 3
3 3 1 3
8 3 0 3 0 3 1 3 3
7 3 0 0 3 0 1 0
3 3 3 2
8 3 0 3 1 3 3 3 2
5 3 0 1 0 0
6 3 0 2 3 0 0
10 3 0 1 2 3 3 0 1 1 3
5 3 1 0 0 3
2 3 3
8 3 3 0 1 2 0 2 3
18 3 0 0 2 1 1 1 1 1 3 3 2 1 3 3 3 3 0
2 3 3
7 3 3 1 3 3 0 3
2 3 3
3 3 0 3
4 3 1 2 0
2 3 3
8 3 0 1 3 3 3 0 2
4 3 1 1 3
10 3 0 3 3 0 2 3 1 2 3
9 3 3 2 1 1 2 0 3 0
21 3 0 3 1 2 1 1 3 2 1 2 0 3 0 1 3 3 1 3 3 0
8 3 0 3 1 0 1 3 3
9 3 1 1 3 0 3 0 1 2
7 3 0 3 1 2 0 3
11 3 0 3 0 1 3 3 0 1 3 3
8 3 3 1 2 3 1 3 0
3 3 3 3
3 3 0 3
2 3 3
14 3 0 3 1 2 1 2 3 2 0 0 2 3 3
13 3 0 3 1 0 1 3 3 0 2 1 3 0
1 3
15 3 3 1 3 0 3 3 3 0 3 1 0 1 3 3
2 3 3
2 3 3
3 3 0 3
5 3 3 0 0 0
8 3 3 0 0 0 3 2 0
19 3 1 1 1 1 1 3 3 3 3 3 3 0 2 3 0 2 0 3
9 3 0 3 0 1 3 3 3 0
14 3 1 1 3 3 0 3 1 0 1 2 1 1 3
4 3 3 3 2
3 3 3 0
10 3 0 3 1 2 3 0 1 1 3
3 3 3 2
7 3 0 3 0 1 2 3
9 3 1 3 1 0 3 2 0 3
7 3 0 3 1 0 1 2
3 3 0 3
1 3
6 3 0 2 3 0 2
6 3 3 0 2 0 3
6 3 0 2 3 0 0
4 3 0 1 0
2 3 3
2 3 1
10 3 0 3 0 1 2 3 0 2 3
3 3 3 2
4 3 3 0 1
11 3 0 2 3 0 1 2 0 3 3 0
7 3 3 0 2 1 3 3
8 3 0 3 0 3 2 0 3
4 3 0 3 0
7 3 0 3 0 3 1 1
2 3 3
16 3 0 3 1 3 3 0 1 2 0 3 1 2 0 3 1
4 3 1 1 3
12 3 0 3 1 2 2 0 0 0 3 0 0
3 3 3 0
4 3 0 3 3
6 3 0 3 1 2 3
2 3 3
17 3 0 3 0 0 2 1 0 1 0 0 1 1 1 2 1 3
1 3
16 3 3 1 3 3 1 3 1 3 1 3 3 3 0 0 0
4 3 0 2 3
2 3 3
2 3 3
10 3 0 3 0 1 3 3 0 0 3
14 3 0 3 0 1 1 3 1 3 1 3 3 2 3
7 3 0 1 2 0 3 0
5 3 0 3 3 0
4 3 3 0 0
10 3 3 0 1 1 2 3 0 0 3
3 3 1 3
5 3 0 3 3 0
2 3 3
4 3 1 1 2
2 3 3
4 3 1 2 0
1 3
18 3 3 0 2 3 1 3 3 3 0 2 1 3 0 3 3 0 3
10 3 0 3 1 0 2 1 0 3 1
9 3 0 2 3 1 1 1 1 2
7 3 1 3 1 3 3 1
2 3 0
7 3 0 3 0 1 2 3
2 3 3
6 3 1 1 3 0 3
5 3 0 2 1 3
6 3 3 0 0 3 0
4 3 0 3 0
5 3 0 3 1 3
6 3 0 3 0 1 2
2 3 3
7 3 3 1 3 0 0 3
5 3 0 3 3 0
34 3 0 1 1 3 3 3 0 1 0 0 3 3 3 1 2 2 1 3 1 3 3 0 2 1 1 1 1 3 1 1 1 3 0
1 3
11 3 0 3 0 1 3 3 1 3 0 0
4 3 0 3 3
5 3 0 3 1 0
5 3 0 3 1 3
9 3 0 2 3 1 3 3 0 2
3 3 3 0
5 3 1 3 0 0
9 3 0 1 3 3 1 1 3 3
1 3
1 3
3 3 3 0
1 3
4 3 0 3 3
20 3 3 1 3 3 3 1 3 3 0 3 0 3 1 3 1 1 1 1 1
8 3 1 3 3 1 2 0 3
17 3 0 3 1 3 0 1 2 2 1 3 0 2 0 3 1 3
2 3 3
10 3 1 3 0 2 1 0 1 3 0
6 3 0 3 0 3 0
5 3 0 3 0 2
4 3 1 1 3
2 3 3
2 3 3
4 3 0 2 3
4 3 1 3 0
8 3 1 0 0 1 1 0 0
6 3 3 0 2 0 3
3 3 0 3
5 3 0 3 0 3
3 3 0 3
8 3 0 3 0 3 0 0 3
9 3 3 2 0 2 3 1 3 3
1 3
3 3 0 3
8 3 3 2 2 2 3 0 2
4 3 0 2 1
3 3 1 3
7 3 1 3 0 0 1 3
8 3 0 3 1 2 0 3 0
3 3 1 3
2 3 3
2 3 3
5 3 1 0 1 3
12 3 3 1 3 3 3 0 1 1 1 1 3
3 3 1 1
7 3 0 3 0 3 0 3
13 3 0 3 0 0 3 1 2 2 0 3 0 3
5 3 3 0 1 0
6 3 0 3 3 0 2
7 3 0 3 0 3 0 0
5 3 0 3 3 0
14 3 0 3 1 0 2 3 0 3 0 1 3 3 0
10 3 0 2 3 0 1 1 1 2 3
4 3 0 3 3
6 3 0 2 1 1 3
4 3 3 0 2
7 3 1 3 0 2 1 3
2 3 3
8 3 3 0 3 3 3 0 0
7 3 3 0 2 0 3 0
10 3 0 3 1 0 1 2 3 1 3
3 3 3 3
2 3 3
4 3 3 2 0
6 3 0 3 0 2 0
24 3 3 1 3 3 0 3 0 1 3 3 0 3 1 3 3 0 0 0 1 0 1 0 2
6 3 2 0 1 3 0
2 3 3
3 3 3 0
9 3 3 1 3 3 0 2 0 0
20 3 1 3 0 2 0 3 1 3 0 3 1 2 2 0 2 3 3 1 3
3 3 3 0
14 3 3 2 3 3 2 0 1 2 2 1 3 0 3
3 3 3 2
5 3 0 3 0 2
3 3 3 0
14 3 1 3 0 3 3 3 3 1 3 3 1 1 1
4 3 3 3 0
8 3 0 3 1 3 0 3 0
2 3 3
8 3 1 0 1 3 1 0 0
3 3 1 3
1 3
2 3 0
12 3 0 3 0 2 3 2 0 3 0 0 3
4 3 1 1 3
3 3 0 3
8 3 1 3 0 1 2 3 3
3 3 0 3
7 3 0 3 0 1 2 1
3 3 0 3
16 3 0 3 1 2 1 2 3 2 0 1 2 3 0 1 2
3 3 1 3
1 3
2 3 0
5 3 0 3 0 0
13 3 3 2 0 2 2 0 3 1 0 2 1 1
4 3 2 0 3
3 3 0 3
3 3 1 3
11 3 1 1 3 0 2 3 1 3 3 0
4 3 3 0 2
11 3 3 1 3 0 3 0 2 3 0 2
19 3 1 1 3 0 0 1 3 1 3 2 2 2 3 1 2 1 1 3
9 3 0 3 1 0 1 3 3 3
3 3 1 3
5 3 0 2 3 0
14 3 0 3 1 0 1 3 3 3 1 3 1 3 0
4 3 1 1 1
2 3 3
1 3
8 3 2 0 3 0 1 1 3
5 3 1 3 0 2
3 3 0 1
9 3 1 2 1 3 3 1 2 0
4 3 0 1 2
3 3 3 0
5 3 0 3 0 1
17 3 0 3 1 3 3 1 3 3 0 3 0 1 3 3 0 3
7 3 3 0 0 0 1 0
2 3 3
4 3 0 3 3
8 3 2 0 3 0 2 1 1
4 3 3 0 2
2 3 3
4 3 0 3 1
15 3 0 3 0 1 3 1 3 1 3 1 1 2 3 3
6 3 3 1 3 2 2
1 3
3 3 1 3
1 3
16 3 3 1 3 3 3 0 3 0 1 3 3 1 0 1 3
19 3 0 2 3 0 2 0 1 3 3 0 3 1 0 1 3 3 3 3
4 3 0 2 3
11 3 1 3 0 0 3 3 1 3 3 3
4 3 3 2 3
6 3 0 3 3 0 2
2 3 0
2 3 3
10 3 0 3 3 2 0 3 1 2 0
17 3 3 1 3 3 0 1 0 1 2 1 2 0 3 1 0 2
5 3 1 3 1 3
6 3 3 0 1 2 1
3 3 0 3
9 3 0 3 3 0 0 1 3 0
2 3 3
5 3 0 3 0 3
1 3
3 3 1 3
10 3 1 2 2 0 3 1 3 3 0
3 3 3 2
5 3 0 3 1 3
10 3 0 3 0 2 0 1 2 1 3
15 3 0 1 3 3 1 2 1 1 1 2 3 2 3 1
8 3 3 0 0 3 0 0 0
3 3 1 3
8 3 0 3 0 3 3 0 0
9 3 3 1 1 3 0 0 1 3
7 3 3 0 2 3 3 0
15 3 1 3 1 3 3 0 1 3 3 3 0 1 1 3
41 3 3 2 3 2 1 1 0 1 2 2 0 3 1 0 1 2 1 3 2 0 3 0 2 3 0 2 0 1 3 3 3 1 3 3 0 3 0 1 0 3
4 3 0 3 3
3 3 1 3
3 3 3 0
3 3 1 3
2 3 3
11 3 1 3 1 3 3 0 1 3 3 3
5 3 1 0 1 3
8 3 0 2 3 0 2 1 3
1 3
5 3 3 1 3 2
1 3
2 3 3
11 3 1 0 3 3 3 2 1 0 2 0
3 3 3 2
7 3 0 3 3 1 3 3
5 3 3 0 1 1
2 3 3
13 3 0 3 0 1 3 3 0 2 3 1 3 3
3 3 3 0
10 3 3 0 0 0 3 3 3 3 0
10 3 3 0 1 1 1 2 0 3 1
10 3 0 1 3 3 1 1 3 0 2
3 3 0 3
2 3 2
9 3 3 0 1 2 3 0 2 0
2 3 1
9 3 3 0 0 1 3 1 1 3
5 3 0 3 0 3
3 3 1 3
2 3 1
12 3 0 1 3 3 3 2 3 1 1 3 3
2 3 0
7 3 3 1 3 3 1 3
4 3 0 2 3
5 3 0 3 1 3
14 3 1 3 1 3 1 3 3 0 3 1 3 0 3
2 3 3
6 3 3 0 2 1 1
2 3 3
6 3 0 2 3 0 1
6 3 3 1 3 3 3
5 3 3 1 3 3
7 3 1 1 3 1 3 3
10 3 3 0 2 0 2 3 0 0 0
10 3 3 1 3 3 0 3 3 3 0
7 3 1 1 1 3 1 3
12 3 3 1 2 3 3 3 1 3 3 3 2
2 3 3
7 3 0 3 3 3 1 3
1 3
4 3 0 3 0
20 3 3 1 3 3 3 1 3 1 3 3 0 1 3 3 0 1 3 3 3
4 3 3 0 1
4 3 1 2 0
9 3 3 1 3 0 1 1 3 1
7 3 1 3 2 0 2 3
2 3 3
11 3 0 1 1 2 3 0 0 1 3 0
2 3 0
12 3 3 1 0 2 0 0 2 2 2 1 3
49 3 3 0 0 1 3 0 2 0 1 3 3 0 3 0 1 3 3 0 1 3 3 3 0 2 0 3 1 0 0 1 3 3 3 0 2 3 1 2 1 1 0 1 3 3 1 0 3 3
4 3 0 3 3
2 3 3
1 3
5 3 3 1 0 2
5 3 0 3 0 3
1 3
2 3 1
2 3 3
3 3 3 2
5 3 0 3 3 3
9 3 1 3 0 1 2 3 1 0
6 3 0 2 2 0 3
4 3 3 0 2
2 3 3
33 3 0 1 3 3 1 3 1 3 3 1 2 2 0 3 1 2 3 0 2 0 3 1 3 0 1 3 2 3 1 3 3 0
1 3
7 3 3 1 3 1 1 3
4 3 3 0 3
2 3 3
1 3
26 3 0 3 1 0 1 2 2 3 1 3 3 0 1 3 3 0 3 3 1 3 3 3 0 0 3
4 3 0 2 3
3 3 0 3
9 3 0 2 3 0 2 1 2 0
5 3 2 0 3 0
6 3 1 3 1 3 3
14 3 0 3 3 2 2 0 3 0 2 2 0 1 3
5 3 0 2 0 0
7 3 3 1 3 3 1 3
1 3
8 3 3 0 0 3 3 0 3
4 3 3 0 2
8 3 0 3 3 1 3 3 3
3 3 3 3
2 3 3
3 3 3 0
5 3 0 3 3 3
25 3 0 3 0 1 1 3 2 2 0 3 0 1 3 2 0 1 3 1 1 1 2 2 0 3
3 3 0 3
8 3 0 2 3 0 2 0 3
3 3 0 3
14 3 0 3 0 3 1 2 1 1 2 3 1 0 0
1 3
9 3 0 3 0 1 2 2 1 3
17 3 3 1 3 3 3 1 2 0 3 0 2 0 3 1 2 3
5 3 1 3 1 0
10 3 3 1 3 2 3 3 3 3 0
7 3 1 3 0 1 0 1
12 3 3 0 1 2 2 0 1 2 3 1 1
5 3 0 3 1 2
1 3
4 3 3 0 2
9 3 1 0 3 3 1 2 1 2
2 3 3
4 3 3 3 0
4 3 1 1 3
2 3 3
13 3 0 3 1 2 2 0 3 1 2 0 0 0
5 3 0 3 3 2
29 3 3 2 0 2 3 2 1 1 2 2 0 3 1 2 1 1 1 1 0 1 2 1 3 1 3 3 0 3
5 3 3 0 0 0
2 3 3
17 3 0 3 0 0 1 3 3 0 3 0 1 3 3 1 0 2
3 3 3 0
2 3 3
5 3 0 3 1 3
15 3 0 3 0 2 1 0 1 2 0 3 1 3 3 0
15 3 3 0 0 1 3 0 0 1 3 0 1 2 3 0
19 3 3 1 0 1 3 3 0 2 1 3 0 1 3 1 3 3 3 3
3 3 1 3
8 3 0 2 3 0 0 0 1
9 3 0 3 0 3 1 3 1 3
1 3
3 3 3 0
6 3 0 3 1 2 3
2 3 0
4 3 1 1 3
4 3 1 3 0
21 3 3 3 0 1 3 3 3 0 2 1 1 3 0 1 2 0 3 3 0 0
8 3 3 1 3 3 3 2 0
2 3 3
2 3 3
9 3 0 3 0 0 3 0 1 2
4 3 0 3 0
2 3 1
20 3 0 1 0 0 3 3 3 1 2 0 0 1 3 0 1 1 1 1 3
8 3 0 3 0 1 3 3 3
3 3 0 1
8 3 3 1 3 3 1 2 1
13 3 0 3 3 0 0 0 3 3 3 0 1 2
9 3 0 3 0 1 0 2 0 3
12 3 3 3 0 1 1 1 2 0 3 1 3
5 3 1 1 0 3
4 3 1 3 0
9 3 0 2 3 1 0 3 3 1
3 3 3 3
4 3 0 2 3
3 3 3 2
6 3 3 0 2 3 3
13 3 0 3 3 0 1 3 1 1 2 3 0 1
4 3 0 3 3
4 3 0 1 0
4 3 1 3 1
9 3 0 3 1 3 0 3 0 2
3 3 0 3
4 3 2 0 3
7 3 3 0 2 1 3 0
8 3 3 1 0 2 1 1 1
3 3 3 0
3 3 3 0
5 3 3 0 0 0
10 3 3 1 3 3 0 2 2 0 3
3 3 0 3
4 3 0 2 3
2 3 3
3 3 3 0
6 3 3 0 2 0 3
2 3 3
2 3 3
4 3 0 2 3
13 3 2 0 3 0 1 2 0 3 3 2 1 0
3 3 1 2
5 3 1 2 3 2
3 3 1 3
12 3 0 3 1 2 3 0 2 0 1 0 3
4 3 0 3 3
4 3 1 3 0
4 3 0 2 3
3 3 0 3
9 3 1 0 0 0 1 3 3 3
4 3 2 0 3
4 3 1 0 0
3 3 0 3
2 3 3
4 3 3 0 2
3 3 0 3
1 3
2 3 3
2 3 3
5 3 3 1 0 3
14 3 3 1 3 3 1 2 1 0 3 2 1 3 0
23 3 0 3 0 2 0 0 0 3 3 1 2 1 2 0 1 1 1 1 1 1 1 1
2 3 3
4 3 3 0 0
4 3 2 0 3
6 3 3 0 0 1 3
11 3 0 3 0 1 3 3 0 3 1 2
9 3 0 3 1 2 2 3 2 0
13 3 0 2 0 0 2 1 1 2 3 0 0 3
7 3 0 3 3 0 3 3
7 3 3 3 0 1 3 1
3 3 0 3
4 3 3 0 1
3 3 3 0
3 3 0 3
2 3 3
10 3 1 1 1 1 1 3 1 3 3
6 3 0 1 3 3 3
2 3 3
5 3 0 3 0 2
11 3 0 3 1 3 1 0 3 3 3 0
1 3
6 3 0 2 3 0 1
6 3 3 0 0 3 0
5 3 0 3 0 3
9 3 3 0 2 0 3 0 2 3
7 3 3 1 3 0 0 1
10 3 0 3 1 2 3 0 2 0 1
17 3 0 3 0 3 1 0 1 3 3 0 0 3 0 1 3 3
2 3 3
1 3
22 3 0 3 0 3 3 1 3 3 0 3 1 2 2 0 3 0 1 0 3 3 0
4 3 3 2 3
17 3 3 0 0 3 3 0 3 0 2 0 3 1 2 1 3 1
4 3 1 2 3
9 3 3 0 2 3 1 3 0 0
4 3 3 0 2
5 3 1 1 3 0
7 3 0 3 0 1 3 3
3 3 3 0
2 3 2
4 3 2 0 3
2 3 0
4 3 3 1 3
2 3 3
1 3
5 3 3 2 1 3
8 3 0 3 0 2 0 0 2
5 3 0 3 0 3
11 3 1 1 3 3 3 1 3 3 0 3
8 3 0 3 1 0 1 2 3
6 3 3 0 0 1 3
12 3 0 3 1 2 0 3 1 3 3 3 0
3 3 1 0
6 3 3 3 1 3 3
13 3 3 3 1 3 3 1 3 3 0 0 1 3
17 3 1 3 1 3 3 1 0 1 3 3 1 2 1 0 1 3
11 3 3 3 0 3 3 0 3 0 1 2
2 3 3
2 3 3
16 3 1 3 3 3 3 1 2 3 3 1 3 3 0 3 3
7 3 0 3 0 1 3 2
6 3 3 1 3 3 3
5 3 1 0 3 3
7 3 3 1 3 3 1 3
11 3 0 3 1 0 1 0 1 3 3 3
23 3 0 3 0 2 0 0 1 3 3 1 3 0 0 0 0 0 0 2 1 3 0 2
16 3 3 2 0 0 2 1 0 3 3 3 1 3 1 3 0
14 3 1 3 1 1 2 0 2 3 1 1 1 1 3
3 3 1 3
12 3 3 0 2 3 1 3 3 3 1 0 0
22 3 0 3 0 1 0 3 1 1 0 1 3 3 3 0 2 2 3 0 1 3 3
3 3 3 2
3 3 1 3
13 3 0 2 3 0 0 1 3 0 0 1 3 1
6 3 3 1 3 3 0
2 3 3
5 3 3 1 2 3
3 3 3 2
14 3 3 0 0 3 3 1 1 1 1 3 0 1 3
10 3 3 0 0 1 3 0 2 0 3
2 3 3
5 3 0 2 3 0
6 3 0 3 1 2 1
1 3
2 3 0
3 3 1 3
6 3 0 3 1 2 1
3 3 1 2
3 3 0 3
9 3 0 3 3 1 3 3 3 0
2 3 0
1 3
1 3
9 3 0 2 2 3 0 0 3 3
2 3 3
4 3 0 3 3
13 3 3 1 3 3 3 3 2 0 0 1 1 3
12 3 0 3 0 2 0 0 2 1 3 3 3
13 3 3 1 3 3 0 3 0 1 3 3 0 2
17 3 0 3 1 1 3 0 1 2 0 3 1 2 1 3 2 1
5 3 0 3 3 0
18 3 0 3 0 1 3 3 3 1 2 3 0 3 0 3 0 2 3
35 3 2 0 1 3 0 2 1 2 1 2 1 1 1 2 1 1 1 0 1 3 3 3 0 1 3 3 3 1 2 2 3 1 3 3
1 3
1 3
7 3 0 1 3 3 0 1
10 3 0 3 3 0 2 0 1 2 3
5 3 0 3 0 1
3 3 3 0
6 3 0 3 0 3 0
2 3 3
7 3 0 3 0 1 3 3
2 3 3
1 3
12 3 0 3 0 3 0 3 3 1 2 0 3
4 3 1 1 3
3 3 3 0
12 3 0 3 3 1 1 2 2 3 1 0 0
2 3 3
15 3 1 3 1 3 3 1 3 3 0 1 1 1 0 1
6 3 3 3 1 1 3
7 3 0 3 0 0 3 0
2 3 3
9 3 0 1 0 2 1 1 1 3
6 3 0 3 1 3 3
2 3 3
10 3 3 2 0 2 1 1 3 1 3
4 3 3 3 0
4 3 0 3 3
1 3
5 3 3 1 3 3
9 3 0 3 1 3 1 2 0 0
9 3 3 1 3 3 1 3 2 0
15 3 3 0 1 1 3 2 0 3 1 3 3 3 0 0
4 3 3 0 0
3 3 3 0
2 3 1
9 3 1 1 3 1 3 3 0 2
3 3 1 3
7 3 0 3 1 2 0 3
2 3 1
11 3 0 3 0 1 3 3 3 1 2 3
5 3 3 0 0 3
7 3 3 2 3 0 1 0
8 3 1 3 0 1 0 3 3
7 3 0 3 3 0 1 1
4 3 0 3 3
6 3 0 3 0 2 3
15 3 3 1 3 3 0 2 3 1 1 1 1 1 1 3
4 3 3 0 0
5 3 0 3 0 3
1 3
4 3 0 3 0
2 3 3
5 3 3 0 2 3
3 3 0 3
37 3 0 1 1 2 3 1 3 3 0 3 1 3 0 3 0 1 2 0 2 0 1 1 1 1 0 1 0 2 1 2 3 1 3 3 3 0
1 3
7 3 1 1 1 3 1 2
5 3 1 1 1 3
9 3 0 3 1 2 2 0 3 0
5 3 3 1 3 3
14 3 1 3 0 2 0 3 1 2 2 0 3 0 2
2 3 3
2 3 1
15 3 1 3 3 1 1 2 3 1 3 3 0 1 3 2
2 3 1
14 3 0 3 3 0 2 1 0 2 3 3 0 2 3
8 3 0 3 3 3 1 2 1
2 3 3
1 3
2 3 3
3 3 1 3
11 3 0 3 1 2 1 2 0 1 2 0
4 3 1 3 1
12 3 3 1 3 3 3 2 3 3 1 3 3
3 3 0 2
22 3 0 3 1 2 2 0 3 0 3 1 2 1 3 0 1 3 3 0 3 1 2
10 3 3 1 3 3 1 2 1 3 0
9 3 3 0 0 1 3 0 1 1
5 3 1 3 0 2
6 3 0 3 0 3 3
2 3 3
3 3 3 2
1 3
18 3 3 0 2 1 1 1 2 0 3 1 0 0 1 3 3 0 1
1 3
7 3 1 3 0 1 1 0
4 3 0 1 1
2 3 3
2 3 3
3 3 1 3
10 3 3 0 0 0 2 3 3 0 2
8 3 0 3 3 1 0 3 1
9 3 0 2 3 1 1 1 1 1
28 3 0 3 1 0 1 0 1 1 3 0 1 2 2 0 3 0 3 0 3 3 0 0 0 0 3 0 3
4 3 0 3 3
11 3 3 1 3 1 1 3 3 2 0 3
8 3 0 3 0 1 1 3 2
4 3 3 1 0
11 3 0 3 0 2 0 0 2 3 3 0
4 3 0 3 0
6 3 0 3 0 2 3
25 3 0 3 0 1 3 3 0 1 3 3 1 1 3 0 3 0 0 3 0 0 1 3 3 3
6 3 0 2 1 3 0
6 3 3 2 1 3 3
3 3 0 3
11 3 3 0 0 1 3 0 0 1 3 0
2 3 3
6 3 3 0 1 1 3
21 3 3 0 1 2 0 3 1 2 2 0 3 1 2 3 1 3 2 1 3 0
2 3 3
1 3
4 3 3 0 2
9 3 0 3 0 1 3 3 3 0
6 3 0 3 1 2 3
3 3 0 3
2 3 3
13 3 1 3 0 1 3 2 2 0 1 3 3 3
10 3 0 3 0 1 1 1 1 1 1
11 3 3 0 1 1 1 1 1 1 1 0
7 3 0 3 1 3 0 2
7 3 0 3 3 3 1 3
13 3 0 2 3 0 2 1 0 3 3 1 2 2
4 3 1 3 0
4 3 0 2 3
29 3 3 1 1 1 1 2 0 1 1 2 0 2 1 3 0 0 0 3 2 3 0 2 3 0 0 3 0 0
2 3 3
17 3 1 3 0 1 2 0 3 0 1 0 1 3 1 0 3 0
10 3 0 3 0 3 1 2 2 0 3
17 3 0 2 3 3 3 3 3 0 1 0 1 2 0 1 1 3
3 3 1 3
2 3 1
4 3 0 3 3
5 3 1 3 0 2
7 3 1 3 0 1 1 0
2 3 3
3 3 0 3
4 3 3 0 0
3 3 3 0
5 3 1 2 1 0
4 3 0 3 0
2 3 3
6 3 3 2 0 1 3
5 3 3 0 1 3
3 3 1 3
2 3 3
15 3 0 3 1 2 0 1 3 1 3 3 1 2 0 2
2 3 3
4 3 0 3 0
23 3 3 1 3 3 1 0 1 2 3 0 0 1 3 1 1 3 2 1 1 2 0 3
4 3 0 3 3
9 3 3 0 1 2 1 1 2 3
6 3 0 3 0 3 0
1 3
3 3 0 3
9 3 0 3 0 3 3 0 0 3
7 3 0 3 3 0 1 1
18 3 0 1 2 0 3 1 0 1 2 3 0 1 2 3 0 3 0
10 3 1 1 3 1 3 0 0 3 3
2 3 0
7 3 3 1 3 0 3 0
11 3 0 3 0 2 0 1 3 0 0 0
2 3 3
5 3 1 3 0 0
9 3 0 3 3 3 1 3 3 0
2 3 0
13 3 0 3 0 3 1 2 0 3 0 0 3 3
8 3 3 0 0 3 0 0 0
3 3 0 3
15 3 1 3 0 2 1 3 0 3 1 0 3 3 3 0
16 3 0 3 0 3 1 2 1 2 3 0 3 2 2 0 3
9 3 3 0 1 3 3 3 0 1
13 3 0 3 0 1 1 3 2 3 1 0 0 3
5 3 2 0 3 0
11 3 0 2 3 0 0 0 1 3 3 3
2 3 3
4 3 1 3 0
3 3 3 2
10 3 3 1 3 3 0 3 1 0 2
2 3 3
14 3 3 1 3 3 3 0 0 1 3 0 0 0 1
24 3 0 3 1 2 2 3 1 3 3 3 1 0 1 1 3 2 1 2 3 1 2 0 3
6 3 0 1 2 0 3
5 3 1 2 0 0
8 3 0 3 1 2 1 1 0
4 3 0 2 3
4 3 3 0 2
5 3 0 2 1 3
6 3 3 0 2 3 3
4 3 3 1 1
7 3 3 1 1 3 0 2
1 3
6 3 3 2 2 2 3
6 3 0 3 1 3 3
1 3
2 3 3
9 3 0 3 0 1 2 1 1 0
1 3
5 3 3 1 0 0
11 3 2 0 3 0 3 1 3 2 0 2
18 3 1 1 3 3 0 2 1 0 3 3 0 3 0 3 0 3 0
5 3 1 3 1 3
5 3 0 2 0 0
9 3 0 1 1 3 3 3 0 3
6 3 3 0 2 3 3
2 3 3
11 3 0 3 1 0 2 2 0 3 0 2
14 3 0 3 1 0 1 2 3 0 1 1 1 3 0
3 3 3 0
2 3 1
1 3
1 3
12 3 3 1 3 3 1 2 2 0 3 0 2
2 3 2
4 3 0 2 3
6 3 0 3 1 2 1
6 3 1 2 0 0 3
3 3 1 3
15 3 1 3 0 3 1 0 1 3 3 3 1 3 3 3
3 3 3 0
11 3 1 3 0 2 0 3 0 1 3 3
2 3 3
3 3 0 3
4 3 2 0 3
4 3 1 3 0
5 3 1 0 1 3
7 3 3 1 2 1 3 0
5 3 0 3 1 0
1 3
6 3 3 1 3 3 0
2 3 3
5 3 1 1 3 0
30 3 1 1 3 1 0 1 1 1 1 1 2 3 1 2 2 3 2 1 1 2 1 3 3 3 0 3 1 1 3
9 3 1 1 1 3 0 1 2 3
3 3 0 3
15 3 0 3 0 3 3 0 2 1 3 2 0 1 0 1
6 3 3 0 2 2 2
4 3 0 3 2
6 3 0 3 2 0 3
16 3 3 2 3 0 2 0 3 1 2 2 0 3 1 2 3
2 3 3
8 3 1 0 3 1 2 0 3
12 3 0 3 1 2 2 3 0 2 1 2 3
17 3 3 1 3 3 3 3 0 0 0 3 0 0 1 1 0 2
4 3 1 1 3
1 3
2 3 0
2 3 0
5 3 1 1 3 3
6 3 3 1 3 3 1
2 3 3
3 3 1 2
2 3 3
10 3 0 3 1 2 3 1 1 1 1
11 3 0 0 3 3 3 0 2 3 0 1
29 3 3 1 3 0 3 1 3 0 3 0 3 0 1 2 2 3 0 2 3 1 3 0 0 0 3 3 3 0
7 3 0 3 3 3 1 0
11 3 3 1 3 3 0 3 1 3 1 3
2 3 0
16 3 1 1 3 3 0 1 2 0 3 0 0 0 3 3 1
8 3 0 3 0 0 3 1 0
10 3 3 0 2 2 0 3 1 1 1
7 3 2 0 3 1 3 3
22 3 3 3 1 1 3 1 3 3 3 0 0 1 3 0 0 3 3 0 1 3 0
6 3 0 3 0 3 0
18 3 0 1 3 3 0 3 0 1 3 3 1 3 0 0 3 3 0
7 3 3 0 2 2 0 3
8 3 0 1 1 3 0 1 0
4 3 0 1 1
3 3 1 2
3 3 3 1
1 3
2 3 3
2 3 3
6 3 1 1 1 1 1
8 3 1 1 3 3 3 3 2
10 3 0 3 0 3 0 3 1 1 3
2 3 3
7 3 3 1 3 3 1 3
3 3 0 3
8 3 0 3 0 3 0 3 3
4 3 0 3 0
2 3 3
12 3 1 1 3 3 1 3 0 3 0 2 0
4 3 0 2 3
3 3 0 3
2 3 3
4 3 1 3 0
13 3 3 0 2 0 2 3 0 0 0 3 0 0
7 3 1 1 1 3 2 3
10 3 0 3 1 0 1 3 3 0 3
15 3 3 3 1 3 3 0 3 0 1 3 3 1 0 2
1 3
3 3 1 3
10 3 3 1 2 1 1 1 1 2 0
8 3 0 3 0 2 3 0 0
13 3 3 0 2 0 3 0 3 1 2 1 0 3
9 3 1 3 1 3 2 0 1 3
6 3 0 3 0 2 1
2 3 3
6 3 0 3 0 2 3
3 3 0 3
1 3
2 3 3
7 3 0 3 0 0 1 0
8 3 3 1 1 0 1 1 2
17 3 0 3 1 2 3 0 2 1 1 1 1 1 3 1 3 0
5 3 0 3 0 3
4 3 1 3 0
5 3 0 3 0 1
6 3 1 1 0 0 1
2 3 3
7 3 0 3 1 0 1 2
7 3 1 3 0 2 3 2
1 3
8 3 1 1 3 3 3 0 1
8 3 3 0 0 1 3 0 2
32 3 3 0 2 3 3 1 1 3 2 1 2 0 3 0 1 2 3 3 1 3 3 3 1 3 3 0 3 0 3 1 3
14 3 0 3 1 0 2 3 3 0 0 3 3 0 0
8 3 1 2 0 2 1 3 0
6 3 0 3 0 2 3
7 3 0 3 0 2 3 0
3 3 3 0
7 3 0 2 3 0 0 3
6 3 0 3 3 0 0
15 3 0 2 3 0 2 1 1 3 3 0 0 3 0 2
2 3 3
8 3 1 1 3 3 1 2 3
6 3 0 3 0 2 1
5 3 3 1 2 3
6 3 0 3 0 2 3
5 3 0 3 0 2
8 3 0 3 1 0 2 0 0
18 3 0 2 3 0 2 0 3 0 1 3 3 0 2 3 1 0 3
6 3 0 1 1 1 3
8 3 0 1 2 2 0 3 3
5 3 3 1 0 2
6 3 3 1 3 3 3
8 3 0 3 0 1 3 3 3
4 3 2 0 3
3 3 3 3
22 3 0 3 0 2 1 1 0 2 0 0 2 1 1 1 3 2 2 0 3 1 3
5 3 3 0 1 1
4 3 3 0 2
5 3 0 3 1 0
4 3 3 0 2
16 3 0 0 2 2 3 1 3 3 0 2 3 0 2 2 2
9 3 0 3 0 3 0 1 3 1
4 3 0 2 3
3 3 0 3
7 3 3 0 1 3 1 2
9 3 3 2 0 0 1 3 0 0
2 3 3
8 3 0 3 1 2 0 3 0
4 3 0 3 3
9 3 0 3 1 2 1 1 0 1
12 3 0 3 0 1 0 1 0 3 1 1 2
1 3
6 3 0 2 1 1 3
2 3 1
13 3 3 2 0 3 0 1 2 3 3 2 0 3
3 3 3 0
12 3 3 1 2 1 1 2 0 3 3 0 0
1 3
10 3 0 3 0 3 0 1 3 2 3
3 3 0 3
6 3 3 0 0 1 3
2 3 3
7 3 0 3 0 1 0 0
2 3 3
2 3 3
1 3
18 3 0 3 0 3 0 2 0 1 0 2 1 2 0 1 2 3 3
6 3 3 1 2 3 0
10 3 2 0 3 0 1 0 1 2 3
7 3 0 3 0 3 1 3
13 3 1 3 0 1 2 0 3 1 3 0 3 3
3 3 0 3
4 3 0 2 3
11 3 1 3 3 1 3 3 1 2 0 3
8 3 0 3 1 3 1 3 0
3 3 0 1
3 3 0 3
23 3 0 3 1 3 0 3 1 2 1 1 1 2 0 3 0 2 2 0 1 3 3 1
3 3 3 0
10 3 3 0 2 0 3 0 1 0 3
1 3
4 3 0 2 3
3 3 2 1
6 3 3 1 3 3 0
7 3 0 3 1 3 3 2
3 3 3 1
2 3 3
2 3 3
5 3 0 2 3 0
8 3 3 0 1 3 3 0 0
5 3 0 3 1 2
2 3 3
4 3 3 3 2
2 3 3
7 3 0 3 0 1 3 3
5 3 3 1 3 2
5 3 1 0 1 3
7 3 3 3 0 3 3 3
10 3 3 1 1 3 2 2 3 1 0
4 3 0 2 3
7 3 0 2 1 3 0 0
3 3 3 2
18 3 1 1 1 3 3 0 1 3 3 0 3 0 1 3 3 0 3
12 3 0 3 1 2 0 3 0 2 2 0 3
52 3 0 3 0 3 0 3 0 3 0 1 3 3 0 3 0 1 3 1 2 0 3 0 2 3 0 2 1 1 3 1 1 1 3 3 2 3 1 3 1 1 3 0 2 1 0 3 0 2 3 0 0
2 3 3
2 3 3
22 3 1 1 3 1 3 3 3 0 0 0 3 3 3 1 2 1 2 0 3 0 1
2 3 3
14 3 0 3 0 3 0 1 2 1 3 1 0 2 2
3 3 3 0
7 3 3 1 3 3 1 2
10 3 0 3 0 3 1 2 3 0 0
11 3 1 3 0 2 1 2 2 0 3 0
1 3
6 3 0 3 1 1 1
5 3 1 3 1 1
4 3 3 3 0
10 3 0 3 0 3 0 1 2 1 1
8 3 3 0 2 1 0 3 3
4 3 1 3 0
6 3 1 3 1 3 0
13 3 3 1 3 3 1 0 1 3 3 0 1 2
6 3 3 3 1 0 2
4 3 1 1 3
15 3 3 0 2 3 1 3 0 2 3 1 2 3 0 0
13 3 1 3 2 0 2 2 0 3 0 2 0 3
28 3 0 3 0 1 3 3 3 1 3 3 1 2 1 3 0 2 3 2 3 0 3 1 2 0 1 1 3
22 3 0 3 1 2 1 2 0 3 1 2 2 3 2 0 3 1 3 2 2 1 3
3 3 3 0
7 3 3 0 2 3 3 0
6 3 1 0 1 3 0
2 3 3
8 3 0 3 1 0 2 0 3
1 3
2 3 3
5 3 1 3 1 3
3 3 0 3
3 3 1 3
5 3 0 3 1 3
5 3 0 3 3 3
2 3 0
10 3 0 3 3 3 3 1 3 1 3
4 3 1 1 3
5 3 0 2 1 3
5 3 0 2 3 0
11 3 1 1 3 3 1 3 1 1 1 3
6 3 0 3 0 0 2
5 3 0 3 1 2
7 3 3 0 0 1 3 0
3 3 3 0
8 3 0 3 0 3 3 3 3
5 3 1 1 3 3
2 3 3
4 3 0 2 3
3 3 0 3
16 3 3 2 0 1 2 1 1 1 0 3 3 0 3 0 2
6 3 3 0 2 1 3
4 3 0 3 0
8 3 3 0 0 3 0 0 2
8 3 3 1 3 0 3 0 3
48 3 0 3 0 1 3 3 3 0 1 3 1 3 1 3 0 1 1 3 1 3 3 3 0 3 0 2 0 1 2 1 1 1 1 3 0 1 3 2 0 1 3 1 3 3 3 0 3
8 3 3 1 1 3 2 1 0
2 3 3
3 3 1 3
22 3 0 3 1 0 1 2 1 1 3 1 3 3 3 1 2 1 1 3 3 1 3
6 3 0 1 0 3 0
1 3
8 3 0 3 1 0 1 1 1
41 3 1 3 0 3 3 3 1 1 1 1 3 1 3 0 0 0 3 3 3 0 3 1 0 2 1 1 1 1 1 2 0 3 0 3 0 1 0 1 2 3
2 3 3
3 3 3 0
15 3 0 3 1 0 1 3 3 0 1 3 3 0 2 3
8 3 0 3 0 2 3 0 0
2 3 3
3 3 1 3
6 3 0 3 2 0 3
2 3 0
1 3
5 3 0 3 1 2
6 3 0 3 3 3 0
5 3 0 2 0 0
4 3 3 0 0
1 3
2 3 3
10 3 3 0 3 0 1 3 3 0 3
7 3 0 3 1 2 1 1
16 3 0 3 1 0 0 2 1 1 3 1 3 1 3 3 2
7 3 3 0 2 0 3 0
4 3 0 3 3
5 3 3 0 2 2
6 3 3 0 0 1 3
10 3 0 1 2 0 1 0 3 1 0
2 3 3
3 3 3 0
5 3 3 0 2 0
15 3 0 2 3 0 2 3 2 1 1 3 0 3 1 3
10 3 3 1 3 3 1 2 3 0 1
7 3 0 3 1 3 0 3
11 3 0 3 3 0 0 3 3 3 2 1
7 3 3 1 3 3 1 3
19 3 1 1 1 3 1 1 3 2 0 1 1 3 0 0 3 3 0 3
8 3 0 3 0 1 3 3 0
9 3 3 0 0 1 3 0 1 3
6 3 1 3 0 2 2
3 3 3 0
3 3 0 3
6 3 3 1 1 1 1
2 3 3
9 3 0 3 3 2 3 2 0 3
5 3 3 1 3 0
2 3 3
9 3 0 3 1 3 0 2 1 2
3 3 0 3
6 3 3 0 2 0 3
10 3 1 2 2 3 0 2 0 1 2
4 3 3 0 0
4 3 3 0 2
7 3 1 3 0 0 3 0
2 3 3
8 3 0 3 0 1 0 0 0
5 3 1 1 3 3
5 3 3 1 0 3
3 3 3 0
9 3 0 3 1 2 2 1 3 3
2 3 3
8 3 0 2 1 3 0 1 0
7 3 0 1 3 3 1 3
6 3 0 3 1 2 3
24 3 3 2 3 0 2 1 1 3 3 0 3 0 3 1 3 3 1 0 2 3 0 0 3
11 3 3 0 2 0 3 1 3 0 0 3
6 3 1 3 0 1 1
3 3 0 1
2 3 3
13 3 1 3 0 2 2 3 1 3 0 2 3 0
10 3 3 0 2 0 3 0 1 3 2
4 3 1 1 3
3 3 3 0
7 3 0 3 1 3 0 0
6 3 3 0 2 0 3
16 3 1 0 3 0 0 1 1 0 1 1 1 2 1 1 2
19 3 0 3 0 2 0 0 1 0 1 1 3 2 0 3 0 1 1 1
25 3 0 1 3 3 0 1 3 3 0 3 1 3 0 3 1 2 1 1 2 0 2 3 0 2
5 3 0 2 3 0
2 3 3
14 3 3 1 3 3 3 1 0 3 3 3 3 1 2
2 3 0
12 3 3 0 0 1 1 3 0 0 1 3 0
1 3
10 3 3 1 3 3 3 1 3 3 3
3 3 3 0
5 3 0 2 3 0
10 3 1 3 1 3 3 1 2 0 3
4 3 3 0 2
1 3
4 3 3 0 2
5 3 0 3 1 3
2 3 3
5 3 3 1 2 3
11 3 3 0 2 0 3 1 3 0 1 0
3 3 1 2
2 3 3
6 3 3 0 2 1 1
2 3 3
2 3 3
5 3 3 0 0 3
5 3 3 1 1 0
6 3 0 3 1 2 3
2 3 0
8 3 3 3 1 3 3 1 2
2 3 3
4 3 3 0 0
5 3 1 3 0 2
3 3 3 0
1 3
3 3 3 2
6 3 1 1 3 0 1
9 3 0 3 0 2 1 0 1 0
5 3 0 1 1 1
3 3 3 0
4 3 3 1 3
11 3 3 0 2 0 3 0 2 0 0 2
3 3 1 3
2 3 3
6 3 1 1 3 3 3
12 3 3 1 3 0 1 2 1 3 2 1 3
2 3 3
6 3 0 3 1 1 3
3 3 0 3
14 3 3 2 0 2 1 2 0 0 1 1 3 1 0
2 3 3
1 3
5 3 3 0 1 1
20 3 0 3 0 1 3 3 1 3 2 0 1 0 1 3 3 3 1 3 0
10 3 0 2 3 1 1 2 3 0 0
10 3 3 2 0 1 1 0 0 1 0
4 3 0 3 0
8 3 2 0 3 0 2 1 2
13 3 3 1 3 3 3 0 1 2 3 1 3 3
5 3 0 3 1 3
2 3 3
1 3
8 3 0 3 0 3 3 3 3
4 3 1 1 3
2 3 3
14 3 3 2 0 0 1 3 0 2 1 3 1 3 3
7 3 2 0 1 3 0 2
5 3 3 3 0 2
14 3 0 1 2 2 1 3 1 3 3 0 1 3 3
2 3 0
8 3 0 3 1 3 3 0 3
19 3 0 3 1 2 1 1 1 1 3 2 0 3 0 2 2 0 3 0
16 3 0 3 1 0 1 3 3 0 3 0 2 0 3 1 3
5 3 1 2 3 2
3 3 0 3
3 3 0 3
6 3 0 1 0 0 1
3 3 1 3
5 3 0 3 0 3
5 3 1 2 0 3
4 3 2 0 3
2 3 3
5 3 0 3 0 3
8 3 3 3 1 3 2 0 3
7 3 0 1 3 3 2 3
5 3 0 2 1 3
8 3 0 3 1 0 1 3 3
8 3 0 3 3 0 0 1 3
7 3 1 3 0 0 1 3
16 3 0 3 1 2 1 1 1 1 0 3 3 1 2 0 3
23 3 3 2 3 0 2 0 3 1 2 2 0 3 0 2 2 2 0 3 0 3 3 0
7 3 3 1 3 3 3 2
10 3 0 3 1 3 0 3 3 3 0
11 3 1 3 0 1 2 0 3 3 3 3
5 3 3 3 0 2
18 3 0 3 0 1 3 3 0 3 0 1 3 2 0 0 2 3 1
8 3 3 3 1 3 3 1 0
3 3 1 3
2 3 3
2 3 3
4 3 1 1 3
2 3 3
2 3 3
3 3 0 3
7 3 0 3 0 1 2 3
10 3 0 3 3 3 0 1 2 1 3
4 3 3 0 0
9 3 3 3 3 1 3 0 1 2
7 3 3 0 2 1 2 3
9 3 3 0 2 0 3 1 2 1
14 3 3 1 2 3 0 3 1 1 3 0 0 1 3
3 3 0 0
3 3 0 3
4 3 0 3 0
6 3 0 3 0 3 3
2 3 3
32 3 3 3 1 3 3 0 3 1 0 1 3 3 0 3 0 0 1 3 3 0 3 0 3 0 3 1 3 1 0 2 1
6 3 0 3 3 2 3
8 3 0 2 1 3 0 1 3
5 3 3 1 3 3
5 3 0 3 0 1
22 3 0 3 0 1 0 0 2 1 2 0 2 0 3 0 3 3 3 0 3 3 3
13 3 1 1 3 3 3 0 1 3 3 3 3 1
3 3 3 0
5 3 0 3 1 3
3 3 1 3
1 3
2 3 3
5 3 0 3 0 2
3 3 0 3
1 3
50 3 3 2 3 0 3 1 0 1 3 3 0 2 0 0 1 3 3 0 3 3 0 2 1 1 3 3 0 2 0 3 3 3 0 3 1 3 0 2 0 3 3 3 1 2 2 1 1 3 0
4 3 0 2 3
6 3 0 3 0 0 3
6 3 3 1 3 3 3
6 3 0 0 3 0 0
5 3 3 0 1 0
5 3 2 2 0 2
3 3 3 1
2 3 2
3 3 0 3
18 3 3 0 2 0 3 0 3 0 1 3 3 3 1 3 3 0 3
3 3 0 1
3 3 1 3
7 3 0 3 3 1 3 3
4 3 3 0 0
3 3 3 2
3 3 1 3
2 3 3
5 3 3 0 2 1
9 3 0 1 3 3 0 1 2 3
24 3 3 3 3 3 1 3 0 3 0 2 0 1 2 1 2 0 3 0 3 0 2 0 3
4 3 2 0 3
2 3 3
23 3 0 3 0 2 3 3 1 1 3 0 2 1 3 1 2 3 0 3 3 0 0 0
2 3 3
28 3 3 1 3 3 1 0 3 3 0 3 3 1 3 0 1 3 3 0 3 3 0 1 2 0 3 1 0
3 3 0 3
12 3 0 3 0 1 2 2 3 2 3 0 2
4 3 0 2 2
2 3 3
11 3 3 1 2 0 3 1 3 3 0 3
1 3
2 3 3
7 3 0 3 0 2 3 0
2 3 3
4 3 0 1 2
4 3 3 0 2
10 3 2 3 0 2 1 0 1 1 1
1 3
11 3 0 3 0 3 0 3 0 1 3 3
6 3 0 3 0 2 2
3 3 1 3
6 3 0 3 0 0 3
3 3 0 3
6 3 0 3 0 2 3
7 3 0 3 1 0 2 3
20 3 0 3 3 0 0 1 3 1 1 1 0 0 1 3 3 3 3 2 0
6 3 0 3 0 2 3
3 3 3 0
6 3 3 1 1 1 3
3 3 1 3
19 3 3 0 2 0 3 1 2 0 3 0 1 1 1 1 0 2 0 3
2 3 3
26 3 0 3 0 1 3 3 0 1 3 3 1 3 0 0 1 3 0 1 1 2 0 3 1 2 3
10 3 0 3 1 0 1 3 3 1 3
4 3 1 1 3
2 3 3
5 3 1 3 0 0
9 3 3 1 2 1 2 1 3 0
3 3 0 3
5 3 0 3 1 0
8 3 0 2 3 1 3 1 3
5 3 1 3 0 1
5 3 2 0 3 0
5 3 0 1 0 0
7 3 1 3 0 2 0 3
7 3 3 0 2 2 0 3
9 3 0 3 0 2 0 3 1 3
12 3 3 2 0 0 3 3 1 0 1 3 3
4 3 3 1 0
7 3 0 2 3 0 0 0
9 3 3 1 3 0 2 1 1 3
1 3
9 3 3 1 3 3 0 3 1 3
8 3 1 3 1 3 1 2 1
3 3 1 3
4 3 0 1 2
16 3 0 3 0 1 3 3 1 2 0 0 3 3 0 3 0
17 3 0 2 3 1 1 0 3 3 0 2 3 0 0 0 1 1
2 3 3
7 3 3 0 2 0 3 0
5 3 0 1 2 1
9 3 1 1 1 1 1 3 1 3
8 3 3 1 3 3 0 2 0
14 3 3 1 3 3 0 0 3 1 2 1 2 0 3
1 3
3 3 0 3
10 3 0 3 0 3 1 3 1 1 1
2 3 3
11 3 3 0 2 0 2 3 3 1 3 0
1 3
5 3 1 3 0 2
11 3 0 1 3 3 1 2 1 1 3 1
5 3 0 3 3 0
18 3 3 1 3 3 0 3 0 1 3 3 0 1 2 1 1 1 0
1 3
12 3 3 1 3 3 2 0 3 0 2 1 2
3 3 1 3
16 3 0 3 0 1 1 3 2 0 3 1 3 3 1 3 0
3 3 1 3
3 3 2 2
15 3 0 2 1 3 0 0 1 3 0 0 0 3 0 0
14 3 0 3 1 2 0 3 0 0 3 3 0 3 0
12 3 0 3 0 3 1 3 0 1 1 3 0
9 3 3 2 1 1 2 1 1 3
11 3 0 3 0 0 3 1 3 0 2 3
1 3
5 3 1 3 3 3
3 3 0 1
7 3 3 1 1 2 0 3
10 3 0 3 1 2 1 1 2 0 3
4 3 0 3 0
5 3 1 1 3 0
2 3 3
6 3 3 1 0 2 0
2 3 0
3 3 0 3
3 3 0 3
3 3 0 3
5 3 3 0 2 0
23 3 3 1 2 3 1 3 0 1 0 1 1 0 1 3 3 0 1 3 1 2 0 3
11 3 1 1 3 0 2 0 3 1 2 1
28 3 3 0 2 1 2 0 2 1 3 3 3 0 1 1 2 0 2 3 1 1 1 1 3 1 1 1 3
4 3 3 0 0
6 3 2 0 0 1 3
8 3 0 3 3 0 1 1 0
9 3 3 0 0 3 3 3 3 3
3 3 3 2
4 3 3 0 2
6 3 3 2 3 0 3
2 3 3
4 3 2 0 3
2 3 0
13 3 0 3 0 2 3 1 3 0 3 0 3 0
17 3 3 0 2 0 3 3 1 0 1 2 3 1 2 0 1 3
6 3 2 0 1 3 0
32 3 0 3 0 1 1 3 3 3 3 3 3 0 1 3 1 1 3 3 3 0 2 3 1 3 3 0 3 0 2 0 3
5 3 0 3 0 1
2 3 3
3 3 0 3
6 3 3 0 0 3 3
4 3 1 1 3
9 3 0 2 2 0 1 3 0 0
5 3 0 3 0 2
2 3 1
11 3 3 0 1 0 2 1 3 1 3 1
8 3 0 3 1 2 1 0 3
4 3 3 0 1
6 3 3 0 0 1 3
5 3 0 3 0 1
2 3 2
14 3 3 0 2 3 1 3 3 0 1 3 3 3 2
6 3 3 3 3 3 2
4 3 3 3 0
2 3 3
2 3 3
2 3 0
1 3
5 3 0 2 3 1
3 3 3 0
12 3 3 3 0 3 3 0 1 3 3 3 0
7 3 3 1 3 3 1 3
4 3 1 3 0
2 3 3
2 3 0
31 3 0 3 3 1 0 2 0 3 0 1 1 3 3 1 0 1 3 3 0 3 0 1 1 1 1 2 3 3 0 0
8 3 3 2 0 0 0 1 3
3 3 3 0
3 3 0 3
9 3 3 0 2 0 3 0 1 0
2 3 3
10 3 1 3 0 1 1 1 3 1 1
13 3 1 3 0 0 3 3 0 0 3 1 2 3
11 3 0 1 0 3 3 0 2 2 2 3
3 3 1 3
13 3 3 1 3 3 3 1 0 0 1 2 1 3
3 3 3 0
12 3 1 0 1 0 0 1 3 3 3 2 2
2 3 3
9 3 3 2 1 1 2 2 3 2
10 3 3 1 3 3 0 1 0 1 0
1 3
4 3 1 3 0
6 3 3 0 1 1 3
7 3 3 2 0 0 2 1
2 3 3
2 3 3
5 3 0 3 1 3
16 3 0 3 0 2 3 0 0 0 1 3 3 3 0 2 3
4 3 1 2 0
3 3 1 3
2 3 0
2 3 3
6 3 3 1 2 3 3
3 3 0 3
1 3
8 3 0 3 1 3 3 0 2
3 3 3 0
7 3 3 1 3 3 3 3
10 3 3 1 3 3 3 1 1 1 3
3 3 3 0
1 3
2 3 3
3 3 1 3
4 3 2 0 3
4 3 0 3 3
2 3 3
10 3 0 2 3 0 1 1 1 1 3
2 3 3
4 3 2 2 0
23 3 3 2 0 1 1 1 2 0 3 0 3 0 3 2 0 3 3 1 3 0 2 3
3 3 1 2
3 3 0 3
5 3 0 3 3 3
8 3 1 1 1 1 1 3 0
7 3 1 1 3 3 0 3
8 3 3 0 2 2 0 3 0
6 3 3 2 0 0 0
12 3 0 3 1 0 1 2 2 3 2 0 3
8 3 0 3 3 3 2 0 0
2 3 3
8 3 0 3 0 3 0 3 0
7 3 1 1 3 3 3 1
16 3 3 2 0 1 2 1 3 0 1 1 3 3 1 3 3
3 3 1 3
10 3 3 2 1 3 3 1 2 3 0
7 3 0 2 3 1 3 3
12 3 3 0 0 3 3 3 2 0 0 1 0
13 3 3 1 3 3 0 0 3 1 2 1 3 0
5 3 3 0 1 3
2 3 0
8 3 3 1 3 3 0 1 2
1 3
1 3
6 3 0 3 0 1 3
5 3 3 0 1 0
11 3 1 0 3 3 3 1 3 0 2 3
5 3 0 3 0 2
10 3 3 2 1 0 1 3 3 0 2
4 3 3 0 1
3 3 1 3
2 3 3
9 3 0 3 1 2 3 1 3 3
11 3 0 3 0 0 0 2 3 1 1 3
4 3 0 3 1
7 3 1 0 0 0 3 3
2 3 1
20 3 0 1 3 3 1 2 0 3 0 2 0 1 3 3 0 2 0 3 0
4 3 0 3 3
5 3 3 1 3 1
2 3 0
8 3 0 2 3 0 0 1 3
6 3 3 0 1 1 0
3 3 1 3
2 3 3
14 3 0 3 0 3 0 0 1 2 3 0 2 3 0
9 3 0 3 3 0 2 0 3 3
2 3 3
6 3 0 3 3 1 1
2 3 3
3 3 3 0
3 3 1 3
2 3 3
3 3 3 0
5 3 3 1 3 2
7 3 0 3 0 0 3 0
4 3 3 0 0
1 3
14 3 3 0 2 1 1 3 3 0 3 1 3 1 3
2 3 0
7 3 1 3 0 0 1 3
2 3 3
29 3 0 3 2 0 0 3 0 1 1 0 2 0 3 0 2 3 0 1 1 2 0 3 0 3 1 3 0 2
3 3 0 1
11 3 3 0 2 0 3 1 2 1 0 1
5 3 2 0 3 0
13 3 3 1 1 1 3 3 2 2 1 1 1 3
9 3 3 0 0 3 3 1 3 3
5 3 1 3 0 2
13 3 0 3 0 3 0 3 0 2 3 0 0 3
11 3 3 0 1 3 0 1 3 3 0 1
7 3 0 3 2 0 3 0
3 3 3 0
8 3 3 1 2 0 1 3 0
6 3 3 0 2 0 3
2 3 3
2 3 3
4 3 3 0 2
2 3 1
18 3 0 2 3 0 1 1 2 0 3 1 0 2 0 2 0 3 3
3 3 0 3
3 3 3 2
3 3 0 3
18 3 3 1 3 2 3 3 3 3 0 1 2 3 0 3 0 1 1
4 3 1 2 0
4 3 3 1 0
10 3 0 3 1 2 3 1 3 3 3
23 3 3 0 0 0 1 0 1 2 0 1 2 3 1 1 1 2 1 3 0 1 1 0
21 3 0 3 0 3 1 3 0 1 1 3 3 3 0 1 0 1 3 1 3 0
3 3 0 3
7 3 0 2 3 0 2 1
7 3 3 1 3 3 0 3
12 3 0 3 0 1 1 0 3 3 1 1 3
2 3 3
4 3 3 0 2
3 3 0 3
10 3 0 2 3 0 2 0 3 0 2
3 3 3 0
8 3 2 0 3 0 0 1 3
41 3 1 1 3 3 3 1 2 1 1 2 0 3 3 0 1 2 0 3 0 1 2 1 0 1 3 3 3 0 1 3 3 0 3 2 0 3 0 0 1 3
3 3 3 2
5 3 1 3 0 0
12 3 0 3 0 1 3 3 0 3 1 2 1
7 3 1 0 3 3 0 3
3 3 3 0
2 3 0
2 3 0
3 3 1 3
6 3 0 1 2 1 3
6 3 1 1 3 3 3
14 3 3 0 2 2 2 3 0 1 0 1 3 3 3
17 3 0 3 1 0 1 3 3 0 3 1 2 3 1 1 3 0
4 3 3 0 2
2 3 3
3 3 3 0
4 3 3 3 2
3 3 1 3
10 3 0 3 1 3 0 3 1 2 3
11 3 1 3 0 1 2 0 3 0 0 3
14 3 2 0 3 0 1 1 2 0 3 3 0 1 0
1 3
1 3
2 3 3
8 3 3 0 1 0 2 1 3
6 3 0 2 1 3 0
2 3 3
30 3 3 2 0 1 1 1 1 1 1 1 1 1 2 3 1 2 3 0 0 0 3 3 3 1 0 1 1 3 0
6 3 1 3 0 1 3
2 3 3
10 3 0 3 0 2 0 1 3 0 3
3 3 0 3
2 3 0
3 3 1 3
6 3 3 1 3 3 3
5 3 3 1 3 1
5 3 0 3 0 3
4 3 3 0 0
10 3 1 3 1 1 1 3 3 3 1
11 3 0 3 3 2 0 1 2 0 2 3
3 3 0 1
1 3
3 3 1 3
6 3 1 3 1 1 3
13 3 1 3 0 2 2 0 3 0 2 0 2 0
7 3 1 3 0 1 2 3
2 3 3
4 3 0 2 3
9 3 1 1 3 0 3 0 2 2
3 3 0 1
4 3 0 3 3
20 3 3 1 3 3 1 2 1 2 3 1 2 1 2 3 1 3 3 0 0
7 3 0 2 3 0 1 0
4 3 0 2 3
5 3 3 1 3 3
2 3 3
6 3 0 3 3 1 2
10 3 0 3 0 1 0 3 3 0 3
6 3 3 0 1 1 3
3 3 1 3
23 3 0 3 1 2 1 1 2 3 2 1 1 0 2 1 1 1 1 0 2 3 2 0
3 3 0 3
17 3 0 3 0 1 3 3 2 0 1 2 0 3 1 2 0 3
11 3 0 3 3 1 3 3 3 1 3 3
2 3 3
7 3 1 3 0 0 1 3
2 3 3
17 3 1 3 3 3 3 1 3 1 1 3 3 3 0 1 0 2
15 3 0 3 0 1 3 3 0 1 3 3 0 3 3 2
8 3 3 2 0 1 1 1 0
1 3
3 3 0 3
5 3 0 3 3 2
17 3 3 1 3 3 1 2 1 1 0 1 2 1 3 0 1 3
2 3 3
4 3 2 0 3
1 3
7 3 0 3 3 2 1 2
2 3 3
6 3 3 0 2 3 2
16 3 0 3 1 2 2 3 1 3 3 0 1 2 1 3 3
14 3 0 3 1 3 1 3 1 1 1 2 1 3 0
4 3 1 1 3
7 3 3 1 2 2 3 2
2 3 3
2 3 3
11 3 3 0 2 3 2 0 0 1 0 0
7 3 0 3 0 1 3 3
5 3 2 0 1 3
13 3 3 1 3 3 0 1 2 0 3 1 2 3
18 3 1 0 3 3 3 1 0 0 2 1 3 1 1 1 1 0 1
7 3 3 0 2 1 0 3
6 3 0 3 1 3 3
9 3 3 1 2 1 1 1 2 3
6 3 3 0 2 0 1
1 3
17 3 3 2 3 1 2 0 2 0 3 1 3 0 3 1 3 3
7 3 1 1 3 3 0 3
2 3 0
3 3 3 0
6 3 3 3 3 0 2
16 3 0 3 1 1 3 3 1 2 1 2 0 3 0 2 3
20 3 0 3 1 2 2 0 3 0 2 0 1 3 3 1 2 1 1 2 2
9 3 0 2 3 0 2 1 3 0
12 3 3 0 2 0 1 3 3 1 1 3 3
4 3 1 1 3
2 3 3
6 3 0 3 2 3 0
15 3 1 3 0 3 3 3 0 0 0 1 1 3 0 1
2 3 3
14 3 1 1 1 1 3 3 0 0 2 0 3 0 2
31 3 3 0 2 3 2 0 1 1 2 3 1 3 3 0 3 1 1 3 0 2 1 1 3 3 2 3 1 3 1 2
4 3 1 3 0
5 3 3 3 0 2
4 3 1 1 1
11 3 0 3 0 1 3 3 1 3 1 3
19 3 3 3 1 3 3 1 3 0 2 0 3 0 2 3 1 1 2 3
17 3 3 2 0 1 3 1 0 0 1 2 3 0 1 3 1 3
8 3 3 1 3 3 0 2 0
2 3 3
19 3 1 1 3 0 1 2 3 0 3 3 0 2 1 1 3 3 1 0
2 3 3
3 3 3 2
12 3 3 0 2 0 3 0 2 3 1 2 3
8 3 0 3 0 1 0 1 0
20 3 0 3 3 3 1 2 1 0 3 0 1 3 3 0 1 3 3 3 2
7 3 1 1 1 1 1 1
3 3 3 0
13 3 3 1 3 0 2 1 3 0 2 1 3 0
2 3 3
2 3 3
5 3 3 1 0 0
2 3 3
29 3 0 2 1 3 3 1 3 3 0 1 0 1 3 0 1 2 0 3 0 1 2 3 3 1 3 2 1 1
2 3 3
5 3 0 3 0 3
4 3 0 3 0
8 3 1 3 1 3 2 0 3
5 3 0 2 1 3
3 3 3 2
4 3 0 3 0
2 3 3
3 3 1 3
1 3
2 3 1
3 3 0 3
8 3 3 0 2 0 3 0 2
3 3 3 0
6 3 3 0 1 1 0
3 3 0 2
11 3 3 0 2 0 3 0 2 0 3 0
2 3 3
3 3 3 0
2 3 3
4 3 1 3 2
6 3 0 3 0 2 3
2 3 3
10 3 0 3 3 0 0 3 3 0 3
10 3 0 3 3 0 1 2 1 3 0
4 3 1 3 0
15 3 1 3 0 2 1 1 3 0 3 3 0 2 0 3
14 3 2 0 3 1 3 3 0 1 3 3 0 2 1
22 3 0 3 1 3 1 0 3 3 1 2 2 0 3 0 1 3 0 1 1 2 3
6 3 3 1 3 1 3
14 3 3 2 3 0 2 0 2 1 1 2 1 3 1
1 3
14 3 0 3 0 2 1 3 0 1 1 3 0 2 2
15 3 0 3 1 1 3 0 1 1 3 2 1 1 0 1
4 3 0 2 3
4 3 3 3 2
6 3 3 1 0 0 3
28 3 3 1 3 3 0 1 2 1 1 3 0 3 0 3 3 3 0 0 1 0 0 1 0 1 2 1 3
2 3 3
6 3 0 3 1 2 3
3 3 1 3
3 3 0 1
7 3 0 3 1 0 1 3
4 3 2 0 3
3 3 3 0
2 3 3
3 3 1 0
10 3 1 3 0 2 0 3 1 3 3
3 3 3 3
3 3 0 1
1 3
7 3 3 2 0 0 0 1
23 3 0 2 3 0 1 2 1 1 3 0 2 3 2 3 0 1 2 0 3 0 3 3
12 3 2 3 1 3 3 0 2 0 2 3 0
4 3 1 1 3
3 3 1 3
4 3 1 3 0
5 3 0 2 1 3
3 3 3 3
2 3 3
11 3 0 3 0 0 1 0 1 3 0 2
9 3 0 3 0 3 0 2 0 3
8 3 3 1 3 3 0 1 1
19 3 3 1 3 3 1 0 2 0 0 2 0 1 0 0 1 2 3 3
10 3 0 1 3 3 3 0 0 0 1
4 3 1 1 3
13 3 0 3 0 2 0 3 0 3 3 3 3 0
4 3 1 3 0
4 3 0 3 0
3 3 0 3
6 3 1 2 1 0 2
10 3 3 0 2 3 1 3 3 0 3
2 3 3
7 3 3 0 2 0 3 3
4 3 3 0 0
7 3 0 3 0 1 3 3
3 3 3 0
6 3 1 1 3 0 3
15 3 3 0 2 1 1 3 0 2 3 0 1 2 0 0
3 3 0 3
12 3 0 3 1 2 1 0 2 1 1 3 3
7 3 3 1 1 1 2 0
3 3 0 1
16 3 1 2 0 0 0 1 1 3 3 1 3 3 0 1 0
3 3 1 3
14 3 3 0 2 0 3 0 0 1 3 3 3 3 3
12 3 0 3 1 2 3 1 3 3 3 0 2
4 3 3 0 2
19 3 1 3 0 2 1 0 3 3 1 3 3 3 0 3 0 1 0 3
7 3 0 3 2 0 3 0
3 3 0 3
18 3 3 0 1 3 3 3 0 1 3 3 0 3 0 3 1 3 3
10 3 3 0 1 2 0 3 3 0 2
9 3 3 0 1 2 3 1 3 3
3 3 3 2
4 3 3 1 1
7 3 1 3 0 2 0 3
16 3 3 2 0 3 0 1 3 3 3 3 1 3 3 3 0
8 3 1 3 0 2 1 0 0
3 3 3 2
7 3 0 1 3 3 3 2
3 3 3 3
7 3 0 3 0 1 3 3
3 3 0 3
4 3 0 2 3
3 3 3 0
4 3 0 1 1
1 3
18 3 1 3 0 2 0 1 0 0 3 3 3 3 0 1 0 3 0
2 3 3
2 3 3
6 3 0 3 0 1 2
7 3 0 2 1 3 1 3
5 3 1 3 2 0
8 3 0 3 0 2 3 0 3
4 3 0 3 3
2 3 0
8 3 1 2 0 2 1 1 3
4 3 1 3 0
21 3 0 3 1 0 1 3 3 0 3 0 1 3 3 1 0 2 2 3 3 3
23 3 0 0 2 3 0 2 1 3 0 0 1 3 0 1 1 2 3 1 0 2 2 3
25 3 3 0 1 1 1 1 1 1 3 1 2 3 0 2 2 0 3 0 2 0 3 2 0 3
3 3 3 0
4 3 2 0 3
2 3 0
3 3 0 3
2 3 3
8 3 0 3 0 1 3 3 3
3 3 1 2
2 3 0
5 3 1 0 2 1
9 3 3 0 3 3 1 2 0 3
10 3 3 0 0 1 3 0 0 1 3
3 3 1 3
10 3 0 0 1 1 2 0 3 3 0
14 3 3 0 0 1 1 3 1 1 1 1 3 1 3
2 3 3
12 3 0 3 0 1 3 3 0 1 2 0 3
3 3 1 3
5 3 3 0 3 3
11 3 3 1 3 3 0 3 3 1 3 3
5 3 1 3 0 0
5 3 2 0 3 0
3 3 3 1
1 3
6 3 0 3 3 2 3
1 3
15 3 0 3 1 2 0 1 3 0 1 3 1 0 1 1
1 3
11 3 3 1 2 0 3 1 3 3 3 1
14 3 0 0 2 0 1 1 2 0 3 0 1 0 2
7 3 3 1 3 1 3 3
4 3 0 3 0
3 3 3 0
1 3
3 3 1 3
4 3 1 3 0
2 3 3
4 3 3 0 0
1 3
1 3
6 3 3 2 0 0 3
3 3 3 2
4 3 1 3 0
3 3 3 3
1 3
5 3 0 3 3 0
2 3 3
3 3 1 3
9 3 0 3 1 0 1 3 3 3
6 3 0 3 2 0 3
10 3 0 3 1 2 0 2 1 3 0
8 3 1 2 1 3 3 0 0
14 3 0 2 3 0 2 0 3 0 2 0 0 2 2
2 3 3
3 3 0 3
5 3 3 0 3 1
6 3 0 3 1 3 0
9 3 3 0 0 1 3 0 0 0
1 3
4 3 0 2 3
1 3
5 3 0 3 1 3
19 3 0 3 1 3 0 1 1 1 2 0 3 0 3 0 2 3 0 1
3 3 3 0
1 3
1 3
7 3 1 3 1 3 3 3
2 3 3
2 3 3
3 3 0 1
1 3
4 3 3 0 2
3 3 2 2
2 3 3
7 3 1 3 0 0 1 3
4 3 0 2 3
3 3 3 0
6 3 1 0 1 3 1
5 3 3 3 0 2
4 3 2 0 3
1 3
11 3 0 3 0 1 3 3 0 3 0 1
12 3 0 3 0 1 3 3 1 3 0 0 0
12 3 1 3 3 2 3 0 2 1 0 3 3
4 3 2 0 3
20 3 0 2 1 3 1 3 1 3 1 3 3 2 1 3 0 3 0 1 2
9 3 0 3 3 1 2 2 0 3
3 3 3 0
6 3 3 3 0 2 2
3 3 0 3
4 3 0 2 3
4 3 0 3 0
12 3 0 3 3 1 0 3 3 1 3 1 3
9 3 0 3 0 1 2 3 1 3
15 3 0 3 1 3 3 0 2 0 3 1 3 0 1 0
17 3 0 3 1 2 0 0 1 1 3 0 0 3 3 0 0 3
4 3 2 0 3
3 3 1 2
2 3 3
4 3 0 2 0
7 3 0 3 0 1 0 3
2 3 3
3 3 1 3
1 3
3 3 1 3
7 3 0 3 0 3 1 3
16 3 0 3 1 3 3 0 2 1 0 0 3 3 3 0 3
3 3 1 2
9 3 3 0 0 0 2 1 3 3
3 3 3 2
8 3 0 3 0 1 3 3 0
22 3 0 3 0 1 2 2 0 3 1 2 0 1 3 1 3 3 3 1 1 2 0
2 3 3
9 3 0 3 1 0 1 3 3 3
3 3 1 3
15 3 0 3 1 2 2 0 3 3 1 3 3 2 0 3
8 3 3 1 2 3 1 3 0
5 3 3 0 1 1
6 3 0 3 1 2 3
15 3 0 1 0 3 3 0 3 1 3 3 3 1 3 3
4 3 3 0 2
7 3 0 1 2 2 0 3
7 3 0 3 1 3 0 1
19 3 0 3 3 2 1 1 2 1 1 0 1 0 0 1 3 0 2 3
6 3 3 1 3 3 3
3 3 3 1
4 3 3 2 0
7 3 3 1 2 3 3 0
7 3 0 3 1 3 1 3
6 3 3 1 1 3 3
9 3 1 3 1 3 3 1 3 0
12 3 3 1 2 0 3 1 3 3 0 3 3
4 3 3 2 0
8 3 0 3 2 0 1 3 0
23 3 0 3 1 2 1 1 1 0 3 1 3 3 1 3 0 0 1 3 1 1 1 1
8 3 0 3 0 3 0 2 3
4 3 3 2 3
7 3 0 3 1 3 1 3
15 3 1 3 0 2 0 3 0 1 1 3 0 3 1 3
3 3 3 0
16 3 0 3 3 1 3 3 0 1 0 1 3 3 1 3 0
2 3 0
12 3 1 3 1 3 3 1 2 0 1 1 1
33 3 3 1 0 0 1 3 3 3 0 3 0 3 1 2 2 0 3 1 0 2 0 2 0 3 0 1 3 3 0 0 3 0
3 3 3 2
7 3 2 3 1 2 1 0
4 3 0 3 0
3 3 0 3
2 3 3
3 3 1 3
15 3 3 1 3 3 0 3 0 3 0 1 1 0 1 3
3 3 0 3
6 3 0 3 1 0 2
2 3 3
3 3 3 3
6 3 0 0 2 1 3
1 3
8 3 1 1 1 1 1 1 1
5 3 1 3 0 2
5 3 1 3 0 0
5 3 0 3 0 1
4 3 1 3 0
6 3 3 0 1 0 1
4 3 1 1 3
9 3 0 3 1 3 2 0 1 3
2 3 3
11 3 0 3 0 1 3 3 0 1 3 3
4 3 0 3 0
9 3 0 3 0 1 2 2 3 0
4 3 3 0 0
4 3 3 0 0
21 3 0 3 0 3 1 3 0 2 1 1 1 2 0 1 2 3 0 1 0 0
5 3 0 3 3 3
7 3 0 3 0 1 3 3
2 3 3
23 3 0 3 0 1 3 3 3 1 1 1 2 0 1 1 3 0 2 0 3 1 2 3
3 3 0 3
2 3 3
26 3 2 3 1 0 1 3 3 0 2 3 1 1 2 3 3 1 0 2 1 2 1 3 0 3 3
2 3 0
4 3 0 2 3
3 3 3 0
3 3 3 0
2 3 3
8 3 0 2 3 0 1 1 0
8 3 3 1 2 0 3 0 2
6 3 0 3 0 2 3
17 3 0 3 0 1 3 3 1 0 2 0 2 0 3 0 1 2
3 3 0 2
2 3 3
5 3 0 3 0 3
2 3 3
6 3 0 2 3 0 0
3 3 3 2
9 3 0 3 0 1 0 0 0 0
3 3 3 0
13 3 3 2 0 0 1 3 3 0 3 1 2 3
1 3
9 3 0 3 1 1 3 3 2 1
4 3 2 0 3
1 3
4 3 0 1 2
3 3 1 3
1 3
9 3 3 0 1 3 0 1 0 2
4 3 3 0 0
2 3 0
7 3 0 1 1 2 0 1
2 3 3
9 3 0 3 3 1 2 2 0 3
9 3 0 3 0 1 1 3 3 0
4 3 1 3 0
19 3 3 0 2 0 1 2 2 3 1 1 3 0 3 0 3 1 2 3
2 3 3
6 3 1 1 3 3 3
3 3 0 3
7 3 3 0 1 1 2 3
6 3 3 0 2 0 3
13 3 3 1 1 0 3 0 0 1 1 3 0 2
1 3
1 3
14 3 0 3 1 2 1 1 1 2 0 2 3 1 3
3 3 0 3
3 3 0 3
6 3 3 1 1 0 0
2 3 3
4 3 0 2 3
5 3 0 3 1 3
2 3 3
2 3 3
2 3 3
2 3 3
2 3 3
5 3 0 2 3 1
7 3 1 3 0 2 0 3
3 3 3 0
9 3 0 3 1 2 1 2 0 3
4 3 1 1 3
6 3 2 0 1 3 0
3 3 3 1
21 3 1 3 1 3 3 0 3 0 1 1 3 3 1 2 2 0 0 1 1 3
3 3 0 3
1 3
3 3 1 2
7 3 1 1 1 1 3 3
12 3 3 1 3 3 1 1 3 0 1 2 3
3 3 0 3
6 3 3 1 3 3 0
4 3 0 2 0
7 3 1 2 0 1 0 2
6 3 0 1 0 1 3
2 3 3
3 3 3 0
9 3 3 2 0 1 1 2 0 3
11 3 0 2 3 0 3 1 2 1 1 0
9 3 0 3 0 1 3 3 3 0
9 3 1 3 0 3 2 3 3 2
5 3 3 1 3 3
4 3 1 0 0
14 3 3 1 3 3 3 0 2 0 3 1 2 1 3
8 3 0 3 0 1 2 1 0
3 3 0 3
4 3 3 0 2
15 3 0 2 3 1 2 1 1 1 3 3 1 1 1 0
1 3
7 3 3 1 3 3 0 2
8 3 0 3 1 3 3 0 0
6 3 3 1 3 3 3
11 3 0 3 0 1 2 1 3 0 3 2
2 3 0
5 3 3 0 2 1
3 3 1 3
10 3 3 1 1 1 1 1 3 3 3
7 3 0 3 3 0 2 1
3 3 0 3
9 3 3 1 3 3 1 3 0 1
4 3 0 3 0
4 3 1 2 0
3 3 3 0
8 3 1 3 0 2 0 3 0
8 3 3 2 1 1 3 0 2
8 3 0 3 0 2 3 1 3
13 3 0 2 3 0 2 0 2 3 0 0 1 3
29 3 0 3 1 0 1 0 0 1 3 2 3 1 2 1 2 0 1 1 1 3 2 1 1 3 3 3 3 3
6 3 0 3 3 2 0
3 3 3 0
7 3 0 2 0 0 0 3
4 3 2 0 3
14 3 0 3 0 1 3 3 3 3 0 1 1 0 2
2 3 2
8 3 0 3 0 2 2 2 3
9 3 3 0 2 3 3 0 0 0
11 3 1 3 0 0 3 0 0 0 1 3
4 3 1 1 3
17 3 3 1 2 1 1 1 1 1 1 1 2 3 1 2 0 3
3 3 3 0
3 3 3 0
1 3
6 3 3 3 1 3 3
9 3 3 0 2 3 2 3 0 3
3 3 3 0
3 3 1 3
3 3 3 0
4 3 0 3 0
3 3 1 3
1 3
7 3 0 3 1 2 1 3
12 3 0 3 2 2 1 1 0 1 3 3 3
6 3 3 2 3 0 3
4 3 0 3 0
3 3 1 3
2 3 3
13 3 0 3 3 1 3 3 1 2 0 1 0 1
4 3 3 0 0
2 3 0
12 3 3 1 3 3 0 2 3 1 2 0 0
8 3 3 0 1 1 1 1 0
4 3 0 2 3
2 3 3
3 3 0 3
12 3 3 2 3 3 1 3 3 3 0 2 3
7 3 0 3 0 2 1 3
1 3
9 3 0 3 3 3 0 3 0 1
7 3 0 3 0 2 3 0
11 3 0 3 0 3 1 3 3 0 2 2
7 3 0 3 1 2 1 2
8 3 0 1 2 1 1 3 3
9 3 0 3 0 2 1 3 0 0
3 3 3 2
3 3 3 2
8 3 1 3 1 1 3 1 3
6 3 1 3 0 3 0
10 3 0 2 3 0 0 1 1 3 0
1 3
4 3 3 2 3
3 3 0 3
4 3 3 1 2
6 3 0 3 0 3 3
16 3 0 3 0 1 3 3 3 0 1 3 0 1 3 3 3
6 3 0 1 0 3 2
5 3 3 0 0 0
1 3
2 3 3
28 3 1 2 0 2 2 0 3 1 3 3 3 1 3 3 0 1 0 1 3 2 1 0 3 3 2 0 3
6 3 1 0 1 3 0
7 3 0 3 3 0 3 3
17 3 0 3 0 1 1 3 3 3 3 3 3 3 0 0 0 1
2 3 2
5 3 0 1 1 1
6 3 0 3 1 2 3
9 3 0 1 3 3 1 3 3 2
2 3 3
15 3 0 2 2 2 3 1 3 3 0 3 0 1 3 3
5 3 0 3 1 2
2 3 0
4 3 0 3 0
13 3 0 3 0 3 0 3 1 1 3 0 2 0
8 3 0 3 0 1 1 3 3
15 3 3 0 1 2 0 3 1 2 3 0 1 1 2 0
2 3 3
3 3 1 3
1 3
2 3 3
2 3 1
6 3 3 1 2 1 2
7 3 1 1 3 3 3 0
14 3 3 0 1 1 1 1 1 2 0 3 3 0 0
9 3 0 3 1 0 0 1 0 0
26 3 1 1 1 0 2 1 1 1 1 3 3 0 1 3 3 0 1 3 3 0 1 0 2 3 3
15 3 3 0 0 1 3 3 1 3 3 0 1 3 3 0
4 3 1 3 0
6 3 3 0 0 0 2
9 3 0 3 1 2 1 1 0 1
4 3 3 0 0
22 3 0 3 0 3 3 1 3 2 3 0 3 3 0 0 0 1 1 0 1 3 1
2 3 3
4 3 3 2 0
6 3 3 0 2 1 0
2 3 3
4 3 1 3 0
3 3 3 0
3 3 0 1
2 3 3
13 3 0 3 0 1 3 3 0 3 3 0 1 3
3 3 0 0
2 3 0
8 3 0 3 1 2 0 3 0
1 3
7 3 0 3 1 3 1 3
8 3 0 1 2 3 2 0 3
12 3 3 2 3 1 1 3 3 3 1 3 3
5 3 0 3 0 2
5 3 0 1 2 1
11 3 3 0 1 1 0 1 3 2 3 0
7 3 3 1 3 3 0 3
3 3 0 3
4 3 1 0 0
12 3 3 1 3 3 3 1 3 3 3 1 3
7 3 1 3 1 3 3 0
2 3 3
14 3 0 3 1 3 3 0 0 1 3 3 0 0 3
8 3 0 3 0 1 2 0 2
11 3 3 0 2 1 0 3 3 1 3 3
6 3 3 3 2 2 3
11 3 3 1 3 3 3 1 3 3 3 0
20 3 0 3 1 2 1 1 1 0 0 0 3 0 1 0 1 3 1 0 3
6 3 0 3 1 3 0
7 3 0 2 3 0 0 0
18 3 3 0 0 0 1 0 1 3 3 0 3 0 1 3 3 3 0
5 3 0 3 3 0
3 3 1 3
4 3 3 2 0
4 3 2 0 3
3 3 0 3
3 3 1 3
4 3 3 0 2
27 3 3 2 3 0 3 0 1 3 3 0 3 0 0 3 0 1 3 3 0 3 0 1 3 1 0 3
3 3 0 3
10 3 3 1 3 3 0 2 3 0 0
2 3 3
9 3 3 0 1 3 2 0 1 3
12 3 3 1 1 3 1 3 0 0 1 1 3
7 3 0 3 1 0 2 0
4 3 3 0 2
6 3 0 3 3 0 1
4 3 3 1 2
3 3 0 3
6 3 3 0 0 1 3
5 3 0 3 3 0
9 3 1 3 1 3 3 3 0 1
3 3 0 3
2 3 3
3 3 0 3
5 3 0 3 0 2
7 3 3 1 2 3 0 2
12 3 0 3 0 1 2 1 1 3 0 1 0
6 3 0 3 3 2 3
3 3 3 2
4 3 0 2 3
5 3 0 3 3 0
4 3 1 3 0
2 3 3
4 3 3 3 2
14 3 0 3 0 1 2 3 0 3 3 0 2 2 3
3 3 3 0
5 3 0 3 3 3
2 3 0
6 3 0 1 3 3 3
2 3 3
8 3 0 3 0 2 0 0 0
4 3 0 3 3
2 3 0
2 3 3
1 3
2 3 3
2 3 3
6 3 3 0 2 1 2
16 3 0 3 0 1 2 2 0 3 3 0 0 1 3 0 2
9 3 0 3 1 1 3 0 1 0
2 3 3
6 3 3 1 2 1 2
3 3 0 3
27 3 1 1 1 1 1 3 1 3 1 1 3 2 0 3 0 0 1 3 0 0 3 3 1 3 0 1
25 3 0 3 1 2 2 0 3 0 0 3 0 1 3 3 0 3 1 2 1 1 2 3 3 2
2 3 3
1 3
25 3 0 3 0 3 0 2 3 0 1 2 1 2 2 0 3 0 2 0 3 1 3 0 3 0
7 3 3 0 1 1 2 3
15 3 3 0 1 1 1 1 2 0 3 0 3 0 3 0
3 3 3 0
3 3 1 3
5 3 0 3 1 2
1 3
9 3 3 1 3 3 3 1 3 3
5 3 3 1 0 0
10 3 3 1 3 3 3 0 3 3 3
12 3 3 1 3 3 1 3 3 0 0 3 3
3 3 3 2
6 3 0 3 0 1 2
5 3 0 3 0 2
3 3 1 3
7 3 0 3 1 2 3 0
1 3
5 3 3 1 3 3
4 3 0 3 0
8 3 0 2 3 0 2 0 3
2 3 3
9 3 2 0 1 1 3 0 1 3
7 3 1 3 0 2 0 2
8 3 2 0 3 0 2 3 2
2 3 3
6 3 0 1 3 3 3
4 3 3 0 2
6 3 0 3 1 3 0
7 3 3 1 3 3 0 2
8 3 0 3 0 3 1 3 3
13 3 3 0 3 3 0 3 1 3 0 2 3 1
3 3 0 3
3 3 1 3
4 3 3 0 0
7 3 0 3 3 3 0 2
1 3
3 3 1 3
5 3 0 3 0 2
15 3 0 2 3 0 0 0 3 3 3 0 1 3 1 3
6 3 1 1 1 3 0
13 3 1 1 3 3 0 3 3 3 0 3 3 0
24 3 3 2 0 1 1 1 1 2 0 3 3 0 2 1 0 3 3 3 1 3 3 3 0
17 3 0 3 1 2 0 3 0 2 1 1 3 3 1 1 1 1
13 3 0 3 1 3 1 3 0 0 3 3 2 0
3 3 0 3
3 3 3 0
1 3
1 3
2 3 1
1 3
21 3 0 1 0 1 2 0 1 3 0 2 0 3 1 2 1 1 1 1 0 2
3 3 0 3
6 3 1 1 1 1 3
2 3 3
16 3 0 3 1 2 2 0 3 0 1 0 3 3 1 3 3
30 3 1 1 1 3 2 1 0 3 0 0 1 0 2 3 3 1 3 0 2 1 3 3 3 0 3 0 1 3 3
6 3 0 3 3 0 2
4 3 1 2 3
5 3 3 2 1 0
12 3 3 1 3 3 1 3 1 1 3 0 0
7 3 0 3 1 2 3 0
2 3 3
8 3 3 0 3 3 0 3 3
2 3 3
26 3 3 0 2 0 2 1 3 0 1 3 2 2 0 2 3 0 2 1 3 1 3 0 2 3 0
13 3 0 3 0 3 0 3 0 3 0 2 0 3
1 3
23 3 0 3 0 1 0 3 3 0 3 1 3 0 2 0 3 0 1 3 3 0 3 0
5 3 0 2 3 0
6 3 0 3 0 3 0
8 3 3 0 2 1 0 0 0
9 3 0 3 1 0 2 2 3 0
6 3 3 1 3 3 3
6 3 0 3 1 1 3
8 3 0 3 3 0 2 0 3
5 3 1 1 1 1
14 3 1 3 0 3 3 0 0 1 3 3 0 2 2
8 3 0 3 3 1 2 1 3
3 3 0 3
12 3 3 1 1 3 1 3 3 1 3 3 0
4 3 1 3 0
7 3 3 0 1 3 2 1
1 3
2 3 3
10 3 2 1 0 3 0 0 1 3 3
23 3 1 3 0 2 1 1 1 3 0 0 1 1 1 1 2 3 1 3 0 2 3 0
3 3 0 3
2 3 0
7 3 0 3 1 2 2 3
13 3 0 3 0 3 0 1 3 3 3 0 3 3
11 3 0 3 1 0 1 3 3 3 2 0
1 3
5 3 0 2 3 0
8 3 0 3 0 3 0 1 2
2 3 3
2 3 3
3 3 3 2
2 3 3
12 3 1 3 0 0 1 3 1 3 3 0 3
6 3 0 3 0 2 3
6 3 0 3 0 0 3
3 3 1 3
11 3 0 3 0 1 2 2 0 3 3 3
3 3 0 3
7 3 3 0 1 1 1 3
4 3 3 0 0
9 3 3 2 3 0 2 2 0 3
12 3 3 1 3 1 1 3 1 3 3 1 3
2 3 3
3 3 0 3
1 3
12 3 3 2 0 2 0 3 1 3 1 1 3
31 3 3 1 3 3 3 0 1 1 2 0 3 1 2 2 0 2 3 0 2 1 2 0 1 1 3 1 0 1 0 0
16 3 0 3 1 0 3 3 0 3 0 3 1 2 1 3 1
4 3 0 2 3
5 3 3 1 0 0
3 3 1 3
11 3 3 3 0 0 0 1 3 3 0 3
3 3 3 0
22 3 0 2 1 1 3 3 1 3 3 1 3 1 3 3 0 1 0 1 3 3 3
12 3 0 3 0 0 0 3 3 1 0 1 0
10 3 1 3 0 0 1 1 1 3 0
2 3 3
6 3 0 3 0 2 0
1 3
12 3 3 0 1 3 2 3 0 2 2 0 3
14 3 0 3 0 1 2 1 0 1 2 1 1 1 3
4 3 0 3 0
17 3 3 1 3 3 3 0 3 3 3 1 1 3 0 1 3 3
3 3 0 3
2 3 3
5 3 3 1 3 3
3 3 0 3
13 3 3 3 1 1 3 1 3 3 0 3 0 1
6 3 0 3 0 3 1
10 3 3 2 3 0 2 1 0 0 0
3 3 0 3
3 3 0 3
2 3 1
11 3 2 0 3 0 2 0 2 2 3 0
9 3 3 1 3 3 0 2 1 3
6 3 3 0 2 0 3
6 3 2 0 1 3 0
2 3 1
5 3 3 2 3 1
5 3 3 3 0 1
3 3 1 3
6 3 3 3 1 0 0
4 3 0 3 0
3 3 3 0
9 3 0 3 0 2 0 3 1 3
3 3 1 3
6 3 0 3 0 2 3
8 3 0 3 1 0 2 0 0
3 3 0 3
3 3 3 0
4 3 3 2 0
25 3 0 3 1 3 3 1 3 3 1 3 1 1 3 0 0 3 3 3 3 0 2 0 0 0
3 3 0 3
15 3 0 3 3 0 2 3 3 3 3 0 0 1 3 3
13 3 1 1 3 0 2 0 3 3 0 1 0 1
7 3 1 1 3 2 3 1
2 3 3
1 3
6 3 0 3 0 2 3
1 3
5 3 1 3 1 3
3 3 3 0
7 3 3 0 2 2 0 3
2 3 0
2 3 3
4 3 0 3 0
12 3 0 3 1 1 1 1 1 3 1 3 0
1 3
2 3 3
14 3 3 3 2 0 1 1 1 1 0 2 0 3 0
3 3 0 3
3 3 0 3
3 3 0 3
20 3 0 3 1 0 2 1 1 2 3 0 0 0 3 3 1 1 3 1 0
1 3
2 3 3
3 3 3 2
1 3
11 3 0 1 1 3 2 1 1 1 1 0
8 3 0 3 0 1 3 3 3
24 3 3 2 0 1 2 0 3 0 2 0 0 0 3 1 0 1 3 3 1 2 0 3 0
16 3 0 3 1 2 0 3 0 0 1 3 0 1 2 0 3
2 3 3
10 3 0 3 1 2 0 3 0 2 2
4 3 3 3 0
3 3 0 3
6 3 0 1 2 1 3
4 3 0 3 3
4 3 3 0 0
6 3 3 3 0 1 0
1 3
8 3 3 1 3 3 0 3 3
14 3 0 1 3 3 0 1 2 3 0 2 3 1 0
3 3 0 3
4 3 0 3 0
5 3 3 0 0 3
9 3 0 1 3 3 3 0 1 3
10 3 0 1 2 1 1 2 3 0 3
1 3
10 3 3 1 3 3 0 1 3 3 1
1 3
2 3 3
10 3 2 0 3 1 3 0 1 0 3
5 3 0 3 0 2
20 3 3 0 3 3 0 2 0 0 2 3 1 0 1 2 1 2 0 3 3
13 3 3 1 1 1 1 1 1 3 3 2 0 3
3 3 3 0
7 3 3 0 1 1 1 1
1 3
2 3 3
3 3 3 0
9 3 0 3 0 1 1 0 0 0
17 3 0 1 0 2 1 1 2 1 2 0 3 3 1 3 3 3
5 3 1 3 0 2
30 3 0 3 1 2 2 3 3 1 3 0 3 1 1 3 1 3 1 1 3 2 2 3 1 3 3 2 0 0 3
11 3 3 0 2 3 3 0 1 1 1 1
5 3 3 0 0 3
3 3 3 1
3 3 0 3
16 3 0 3 0 2 0 2 3 2 1 1 2 1 3 1 3
1 3
6 3 3 2 0 2 0
20 3 0 3 3 0 1 1 1 1 1 3 2 1 3 1 3 3 3 1 0
9 3 0 1 0 2 0 0 2 0
2 3 3
3 3 3 0
1 3
3 3 0 1
14 3 3 3 1 0 0 2 0 3 1 2 0 1 3
4 3 1 1 1
4 3 0 3 3
3 3 0 3
16 3 3 1 3 3 3 0 3 3 1 0 0 0 2 3 2
2 3 3
2 3 3
12 3 0 1 2 1 1 1 1 3 0 3 0
4 3 3 3 2
7 3 0 3 1 2 3 0
16 3 1 2 0 2 0 3 1 3 3 1 1 3 0 1 3
2 3 0
4 3 0 2 3
5 3 0 3 1 2
5 3 0 3 1 0
4 3 3 0 0
11 3 1 1 1 1 1 1 1 3 3 3
2 3 3
6 3 1 3 1 1 1
5 3 0 2 3 0
4 3 0 3 0
6 3 0 3 1 1 3
2 3 0
2 3 3
18 3 3 3 0 1 2 0 3 0 1 2 3 2 0 0 0 1 3
3 3 1 3
7 3 0 3 3 1 3 3
9 3 1 3 0 1 1 1 1 1
2 3 3
7 3 1 3 1 3 3 3
4 3 3 0 0
23 3 0 2 3 0 0 3 0 0 0 3 3 1 1 2 3 0 0 1 1 3 3 0
15 3 0 3 1 0 2 1 0 1 0 1 3 3 0 2
1 3
21 3 3 1 3 3 3 3 0 2 0 2 2 2 1 3 0 2 2 0 3 0
3 3 0 3
2 3 3
13 3 3 0 1 0 2 0 3 3 0 1 1 1
13 3 3 0 0 1 3 0 1 1 2 0 2 3
5 3 2 0 1 3
1 3
2 3 3
2 3 3
8 3 0 3 1 3 0 2 1
1 3
3 3 3 3
4 3 3 3 0
2 3 0
11 3 3 0 2 1 1 3 3 0 2 3
6 3 1 3 1 2 3
6 3 3 1 0 3 1
8 3 2 0 3 0 0 3 3
27 3 0 3 1 0 2 1 1 3 3 0 2 2 0 3 1 1 1 1 1 3 1 1 2 3 1 0
4 3 0 1 0
16 3 1 1 3 3 1 3 0 2 0 1 1 3 1 1 3
3 3 1 0
3 3 0 1
2 3 3
4 3 1 1 3
14 3 0 3 1 0 2 3 1 1 2 3 0 3 3
10 3 0 3 1 1 3 1 3 0 0
7 3 3 1 3 3 0 3
14 3 1 3 0 1 2 0 3 1 3 3 0 2 1
13 3 0 3 0 2 0 0 1 3 3 1 3 3
10 3 3 1 3 3 0 3 3 3 3
3 3 3 0
20 3 1 3 1 1 1 3 0 1 1 2 0 3 1 2 0 3 0 0 3
5 3 0 3 3 2
2 3 3
6 3 0 3 1 3 3
5 3 1 3 0 0
10 3 3 0 1 1 3 2 1 2 0
18 3 0 1 3 3 3 0 3 3 3 1 3 3 0 1 2 3 0
18 3 0 2 3 0 2 3 2 0 2 0 1 3 3 3 1 3 3
15 3 3 1 1 3 0 3 0 3 0 3 2 1 3 0
3 3 0 3
8 3 1 1 3 0 2 1 3
2 3 3
11 3 1 1 1 1 1 1 3 1 1 3
1 3
3 3 1 3
1 3
8 3 0 3 0 1 3 3 0
7 3 1 2 3 3 1 3
8 3 3 0 1 0 0 0 3
5 3 1 1 3 3
2 3 1
9 3 1 2 0 2 0 2 1 3
7 3 3 0 2 0 3 3
9 3 1 1 3 3 0 2 3 0
9 3 3 1 3 3 3 0 3 0
1 3
3 3 3 0
1 3
4 3 0 3 3
17 3 0 0 1 1 0 2 0 3 1 2 1 1 1 1 1 0
6 3 2 0 3 0 2
2 3 3
12 3 3 1 2 1 1 0 2 3 0 3 0
3 3 3 2
10 3 3 2 0 2 1 1 1 2 0
6 3 0 3 0 3 3
6 3 3 0 2 3 2
2 3 3
12 3 0 3 1 2 0 1 0 2 1 3 0
13 3 0 3 1 3 0 3 3 2 0 1 2 3
1 3
5 3 3 2 3 2
2 3 3
10 3 0 3 0 3 0 1 3 3 1
5 3 2 0 0 3
18 3 0 3 1 3 0 2 0 1 0 3 3 1 2 2 0 3 0
15 3 3 0 2 3 3 0 2 0 2 1 3 1 3 0
2 3 0
13 3 3 0 1 1 0 1 1 1 2 1 1 0
12 3 0 3 0 1 2 1 3 0 1 1 2
6 3 3 1 3 1 2
12 3 0 3 1 3 0 3 1 0 1 3 3
6 3 3 1 3 3 3
2 3 3
26 3 3 1 3 3 0 3 1 2 1 0 2 0 3 3 1 3 3 3 0 3 0 1 3 3 0
28 3 0 1 2 0 3 1 3 3 0 1 2 1 2 0 3 1 0 3 3 0 3 1 2 1 1 3 1
7 3 0 3 1 2 0 3
6 3 3 1 3 3 0
6 3 3 1 3 3 2
12 3 0 3 0 2 3 1 1 1 1 2 3
4 3 1 1 3
15 3 2 0 0 1 1 3 0 1 2 0 0 0 0 3
9 3 1 1 1 3 0 1 1 3
2 3 0
13 3 1 3 1 3 0 0 0 2 0 0 0 3
5 3 3 3 0 2
5 3 0 2 1 3
2 3 3
13 3 0 3 1 3 1 3 1 3 3 3 2 0
3 3 3 2
14 3 2 0 3 0 2 0 3 0 1 3 3 1 3
17 3 0 1 2 0 3 0 1 2 1 3 3 1 3 1 0 3
3 3 1 1
4 3 0 3 0
17 3 0 3 0 2 3 1 0 3 3 0 3 1 2 2 0 3
6 3 1 1 3 3 0
2 3 3
3 3 3 0
7 3 3 1 3 3 1 3
5 3 2 0 3 0
3 3 0 3
4 3 3 0 0
3 3 0 3
4 3 1 2 0
13 3 0 2 1 3 1 2 3 0 3 1 2 3
15 3 1 3 1 0 3 0 2 0 0 2 0 1 2 3
12 3 0 3 1 2 0 3 0 2 2 0 3
2 3 1
13 3 0 3 1 3 3 1 1 1 3 0 3 3
5 3 3 1 3 3
6 3 1 3 0 1 3
39 3 0 3 0 1 3 3 0 3 1 2 1 3 3 3 1 0 3 3 0 3 2 1 1 1 2 3 1 3 3 0 3 0 2 0 0 0 1 3
16 3 0 3 0 3 1 3 1 3 0 2 1 1 3 2 3
21 3 1 1 3 0 3 0 0 3 0 0 3 0 2 1 0 1 0 3 0 3
11 3 1 3 1 3 3 0 2 0 0 2
4 3 0 2 3
2 3 3
30 3 3 1 1 1 3 0 1 1 2 0 2 3 1 3 3 0 3 0 0 1 3 3 2 0 3 0 1 1 0
3 3 0 3
23 3 1 0 1 3 0 1 3 0 0 1 3 3 3 0 1 3 0 3 1 1 1 3
4 3 1 1 3
5 3 3 0 1 3
3 3 1 2
5 3 0 3 3 1
4 3 3 0 0
4 3 0 3 0
2 3 3
18 3 3 0 0 3 3 1 3 3 1 3 2 2 0 1 1 1 3
2 3 3
3 3 1 3
6 3 0 3 3 0 0
4 3 3 0 0
5 3 0 2 3 0
5 3 0 3 1 0
9 3 3 0 2 0 3 0 1 2
6 3 3 0 1 0 1
1 3
5 3 1 1 3 0
3 3 3 0
7 3 0 3 3 1 3 3
3 3 1 2
2 3 3
4 3 0 3 0
17 3 3 1 3 2 2 0 3 1 2 1 2 0 3 0 1 3
11 3 3 3 3 2 0 1 3 0 0 0
3 3 1 3
2 3 3
3 3 3 1
4 3 1 2 2
3 3 0 3
8 3 3 0 1 1 2 0 3
2 3 0
3 3 3 0
12 3 0 3 3 0 2 1 0 3 3 0 3
1 3
5 3 0 2 3 0
9 3 0 3 0 1 2 1 1 1
13 3 3 1 1 3 3 2 2 3 1 3 3 3
19 3 3 0 1 1 2 0 3 1 2 2 3 1 2 3 0 3 0 3
7 3 0 3 1 3 1 3
4 3 0 3 3
9 3 3 0 1 0 0 3 3 0
4 3 0 2 3
8 3 0 3 0 2 2 2 3
15 3 0 3 1 2 0 3 0 1 1 2 3 2 3 2
1 3
11 3 3 2 0 1 0 3 3 0 3 0
4 3 3 1 2
6 3 3 2 2 0 3
6 3 0 3 2 0 3
7 3 3 2 0 2 0 3
2 3 1
5 3 1 3 0 2
8 3 3 1 3 3 3 0 0
3 3 3 0
16 3 0 3 1 3 3 1 1 1 1 1 1 1 3 1 3
9 3 0 3 0 3 1 3 0 3
3 3 1 3
3 3 0 3
26 3 3 1 2 1 0 0 3 1 2 0 1 0 2 3 3 2 0 0 3 0 0 2 2 0 3
8 3 0 3 2 3 0 1 3
8 3 0 3 1 0 1 3 3
3 3 1 3
6 3 0 3 0 3 0
16 3 0 3 1 2 3 0 0 1 3 0 0 0 3 3 3
26 3 0 2 1 1 3 3 3 0 1 3 3 3 0 1 1 1 0 1 1 0 1 1 3 1 0
4 3 1 3 2
11 3 0 3 1 2 1 1 1 1 3 3
1 3
5 3 3 0 0 0
16 3 3 2 1 1 2 2 0 3 1 2 1 1 3 1 2
4 3 0 3 0
21 3 0 2 3 0 2 0 3 0 1 2 2 0 3 1 3 3 0 3 0 3
4 3 0 2 3
7 3 3 0 0 1 3 0
18 3 0 0 2 1 3 3 3 3 1 2 2 1 1 3 0 2 0
6 3 0 3 0 3 3
31 3 3 2 2 2 3 0 2 0 3 0 1 3 2 0 0 2 0 3 1 3 2 3 0 2 1 3 0 0 1 3
3 3 3 2
2 3 1
16 3 0 2 3 1 3 3 0 2 3 1 1 3 3 3 2
2 3 0
19 3 0 3 0 0 3 1 3 1 3 1 3 0 0 3 3 1 1 3
16 3 1 1 3 3 2 0 0 1 2 0 3 0 2 3 2
3 3 0 0
17 3 3 3 1 3 3 0 1 3 3 0 3 0 1 0 1 0
7 3 3 0 2 0 2 3
3 3 0 3
5 3 1 0 3 0
2 3 1
5 3 0 3 0 2
5 3 3 0 0 0
10 3 1 3 0 2 1 1 1 2 3
10 3 3 0 3 3 0 3 0 2 1
3 3 0 3
2 3 3
4 3 0 3 3
32 3 3 2 0 0 3 0 1 3 3 3 2 3 3 0 1 2 0 3 1 3 0 0 2 3 1 3 3 3 0 1 3
4 3 0 2 3
4 3 0 3 0
26 3 1 3 0 2 0 3 0 1 3 3 1 3 3 0 1 1 1 1 1 1 3 3 3 3 3
5 3 3 1 0 3
11 3 0 3 3 0 2 0 1 3 3 0
10 3 0 3 0 1 2 0 3 0 1
13 3 1 3 1 3 3 1 0 1 3 3 0 2
4 3 2 0 3
3 3 1 1
14 3 1 3 0 1 1 2 0 3 0 3 0 1 2
2 3 0
19 3 3 1 3 3 3 0 1 1 2 0 3 1 3 0 0 2 3 1
6 3 0 3 3 2 0
10 3 0 3 0 1 3 3 3 2 0
3 3 1 3
4 3 1 3 2
1 3
9 3 3 1 3 3 1 0 2 3
3 3 0 3
28 3 0 1 2 0 2 3 0 0 3 3 0 1 3 1 3 3 2 0 1 1 3 0 1 2 0 2 3
12 3 0 3 0 1 3 3 1 3 1 3 3
6 3 0 1 2 0 2
12 3 0 3 0 2 3 0 2 3 2 0 3
5 3 0 2 1 3
6 3 3 0 1 1 1
2 3 1
13 3 1 3 0 1 3 2 3 1 0 2 3 0
2 3 3
7 3 1 3 0 0 3 3
8 3 1 1 3 0 1 2 3
4 3 3 2 0
16 3 0 3 3 1 3 3 3 1 2 1 3 0 1 1 3
3 3 0 3
6 3 0 3 1 0 2
3 3 0 3
5 3 0 3 1 0
2 3 1
4 3 3 1 3
3 3 1 3
2 3 3
2 3 3
3 3 3 0
2 3 3
3 3 3 3
1 3
5 3 2 0 3 0
1 3
8 3 0 3 2 0 3 0 2
4 3 2 0 3
8 3 1 1 3 0 0 1 3
3 3 0 3
2 3 3
8 3 0 3 0 1 3 3 3
1 3
9 3 0 3 0 1 3 3 1 3
4 3 3 0 2
3 3 3 2
1 3
3 3 3 3
5 3 1 0 3 3
14 3 0 3 0 1 3 3 0 2 3 2 0 1 3
7 3 0 3 0 0 3 0
8 3 0 3 3 0 0 1 3
5 3 0 3 3 0
3 3 3 0
16 3 3 2 0 3 3 0 2 1 0 3 3 0 2 3 0
13 3 0 3 1 2 1 2 3 0 3 3 3 0
1 3
6 3 0 2 1 1 3
3 3 3 0
4 3 3 2 1
9 3 0 3 0 1 3 3 0 3
18 3 0 3 0 1 3 3 0 2 3 0 3 1 0 1 0 3 1
9 3 2 0 1 3 0 1 0 3
1 3
2 3 3
2 3 3
2 3 3
6 3 0 3 0 1 2
3 3 0 3
14 3 0 3 0 1 1 2 0 0 1 2 0 3 3
13 3 0 3 3 0 0 0 2 1 1 2 2 0
1 3
2 3 0
17 3 3 3 3 2 0 3 1 3 3 0 3 0 3 2 0 3
12 3 0 3 0 3 1 0 1 3 3 0 3
10 3 0 3 0 1 3 3 0 0 3
3 3 0 3
1 3
7 3 0 3 0 1 0 0
10 3 2 0 3 0 2 2 0 3 0
2 3 3
33 3 3 1 0 2 0 3 3 1 3 3 3 0 0 3 3 1 0 1 0 1 2 1 1 1 2 1 3 0 1 2 0 3
3 3 1 1
6 3 3 2 0 0 3
2 3 3
3 3 3 0
4 3 0 3 3
5 3 0 3 0 2
9 3 0 3 0 1 3 3 3 3
3 3 0 1
4 3 0 2 3
4 3 3 0 0
3 3 0 3
3 3 3 3
2 3 3
1 3
2 3 0
14 3 0 3 1 3 3 1 1 1 1 1 3 1 3
14 3 3 1 2 1 3 0 2 1 2 0 0 1 3
2 3 3
5 3 3 0 0 0
28 3 3 1 2 1 3 3 3 0 1 3 3 3 0 2 0 0 2 1 1 1 0 0 3 0 1 3 3
3 3 1 3
12 3 0 3 1 3 0 3 1 3 0 1 0
5 3 0 2 1 3
10 3 0 3 0 1 3 3 3 3 3
13 3 3 0 1 1 3 2 2 0 1 1 1 0
2 3 3
3 3 0 3
4 3 3 2 0
2 3 3
4 3 3 0 0
5 3 2 0 1 3
17 3 3 0 1 1 2 3 1 2 1 1 1 1 2 1 3 0
4 3 3 0 0
2 3 3
3 3 3 0
9 3 0 3 3 1 3 3 3 0
5 3 0 3 0 3
14 3 3 0 2 0 1 2 0 3 1 3 3 1 3
4 3 0 2 3
7 3 0 3 0 1 0 2
6 3 3 0 1 3 1
3 3 1 3
2 3 3
2 3 1
5 3 0 1 2 3
6 3 0 3 0 1 2
5 3 0 3 3 0
3 3 1 3
2 3 3
11 3 3 0 2 0 3 0 3 0 2 3
2 3 3
1 3
12 3 0 3 0 1 3 3 0 3 0 0 2
3 3 0 3
16 3 3 0 2 0 3 0 1 3 3 1 3 0 0 1 3
4 3 3 2 0
4 3 3 2 1
9 3 0 3 0 1 3 3 0 3
3 3 1 1
11 3 0 3 0 2 1 1 2 2 0 3
12 3 3 1 1 3 1 3 3 2 0 0 0
4 3 1 1 3
2 3 3
6 3 3 0 2 1 0
3 3 1 3
6 3 0 2 1 1 3
1 3
2 3 3
3 3 3 3
2 3 3
8 3 0 3 0 1 3 3 3
10 3 0 3 1 2 2 3 1 3 3
2 3 3
11 3 0 0 2 0 0 1 3 3 3 2
4 3 0 2 3
4 3 3 1 0
3 3 0 3
11 3 3 2 0 0 1 3 1 3 3 3
6 3 0 2 3 0 0
3 3 0 3
5 3 2 0 0 3
4 3 3 3 0
3 3 0 3
8 3 0 2 3 0 2 0 3
11 3 3 0 2 0 2 0 3 2 3 3
29 3 0 3 1 2 0 2 0 3 0 1 1 3 1 1 3 0 1 2 0 3 0 2 3 1 1 2 2 3
3 3 3 2
25 3 0 3 1 3 1 1 3 3 3 0 1 3 3 0 3 0 3 3 1 2 1 3 2 3
16 3 3 0 1 2 0 3 1 3 0 3 3 0 2 1 3
7 3 3 1 3 3 3 0
2 3 3
4 3 3 0 1
3 3 0 3
21 3 1 3 1 3 3 1 2 1 3 3 1 2 3 0 2 2 0 3 0 0
5 3 3 1 3 2
2 3 3
2 3 3
5 3 1 1 3 0
3 3 0 3
8 3 3 0 1 2 1 3 0
1 3
7 3 3 1 0 1 3 0
14 3 0 3 0 1 1 3 0 3 3 3 1 2 0
9 3 0 3 1 0 1 2 3 0
5 3 3 1 3 3
12 3 0 3 0 1 3 3 0 2 2 2 3
4 3 0 3 3
8 3 0 3 1 2 0 3 0
6 3 0 3 3 0 0
26 3 3 1 3 3 1 0 3 3 0 1 2 1 1 3 1 1 3 1 1 1 1 3 3 0 3
6 3 0 3 3 2 0
3 3 3 3
9 3 3 0 2 0 3 1 2 3
11 3 3 1 3 0 3 1 2 2 0 3
3 3 1 3
3 3 0 3
8 3 0 3 0 3 1 0 2
7 3 0 3 0 1 3 3
7 3 3 1 3 3 1 2
1 3
2 3 3
8 3 0 3 1 0 2 0 0
2 3 3
10 3 0 3 1 2 2 0 3 1 3
1 3
25 3 0 1 0 1 2 0 3 0 1 2 0 3 3 3 1 0 1 3 3 0 2 3 0 2
12 3 0 3 0 3 0 2 3 0 0 3 3
12 3 0 3 1 3 0 3 3 0 0 1 3
2 3 3
4 3 3 2 0
2 3 3
2 3 0
6 3 0 3 1 2 3
15 3 0 3 0 1 3 3 0 3 3 1 3 3 0 1
9 3 3 3 1 0 0 3 1 3
13 3 0 3 3 3 2 0 3 0 2 0 3 0
2 3 3
7 3 3 0 0 0 1 0
11 3 1 2 3 1 2 3 0 2 0 3
16 3 3 1 0 1 0 0 2 3 1 3 3 3 1 3 3
2 3 3
6 3 3 0 1 1 0
16 3 3 0 2 3 2 0 2 0 3 3 0 1 3 0 2
9 3 3 1 3 3 3 2 3 1
2 3 3
3 3 3 1
2 3 3
25 3 1 3 1 3 0 3 0 3 1 0 1 2 1 2 1 2 0 1 2 1 2 0 3 0
5 3 3 1 3 3
6 3 0 3 1 3 0
3 3 0 2
9 3 0 3 0 3 0 1 3 2
3 3 3 0
4 3 2 0 3
12 3 0 3 0 2 3 1 1 2 0 1 3
3 3 3 0
14 3 3 0 1 1 0 1 2 1 1 2 1 1 3
4 3 3 0 0
7 3 0 3 1 2 0 3
5 3 0 3 0 3
2 3 3
3 3 3 0
11 3 0 3 0 3 0 1 3 3 0 1
6 3 0 3 3 2 1
6 3 0 3 1 3 3
3 3 3 1
4 3 3 0 2
6 3 0 3 1 3 3
35 3 3 3 1 1 1 3 0 3 3 3 1 1 3 3 3 0 1 3 0 1 3 3 1 3 0 0 3 3 3 3 3 0 2 3
10 3 3 1 3 3 0 1 3 3 0
7 3 1 3 0 2 0 3
7 3 3 0 1 1 2 3
1 3
12 3 3 1 3 3 0 3 0 1 3 3 0
3 3 1 0
10 3 1 1 3 0 3 0 1 3 3
14 3 3 0 1 0 1 3 0 1 2 3 0 1 0
6 3 3 0 0 3 3
3 3 1 3
3 3 1 3
2 3 3
1 3
3 3 0 3
1 3
3 3 3 0
3 3 1 3
4 3 3 0 2
8 3 3 1 2 1 1 3 0
6 3 3 1 2 1 1
5 3 3 1 2 3
8 3 0 3 0 1 0 1 2
17 3 0 3 1 0 1 0 0 2 1 1 1 2 0 2 3 3
1 3
4 3 0 3 0
8 3 0 3 1 1 1 1 1
1 3
7 3 3 0 2 2 0 3
6 3 0 3 0 2 0
2 3 3
4 3 1 3 0
3 3 0 3
11 3 0 3 1 3 3 1 3 3 0 1
10 3 0 3 1 2 1 1 3 0 2
32 3 1 3 1 3 3 0 3 0 2 0 1 0 1 3 3 0 3 1 0 1 3 3 1 3 3 0 1 1 1 0 1
20 3 0 3 1 0 1 1 3 0 1 0 3 2 1 3 1 3 3 2 3
2 3 3
7 3 0 3 1 3 0 1
2 3 0
2 3 1
10 3 3 3 2 0 1 2 0 1 3
11 3 1 1 3 0 2 0 3 1 0 2
10 3 3 0 1 2 0 3 3 2 0
20 3 1 0 1 1 2 1 3 0 2 0 1 3 3 0 2 3 1 0 0
1 3
6 3 0 3 1 2 3
9 3 2 0 1 3 1 3 1 3
4 3 1 1 3
5 3 3 1 3 3
8 3 0 3 0 1 2 0 2
11 3 0 3 1 2 1 1 1 3 0 2
2 3 3
17 3 1 1 1 3 2 1 2 3 2 0 1 0 1 3 1 2
2 3 3
16 3 3 1 2 1 1 1 1 2 0 3 1 2 0 3 0
3 3 3 0
9 3 0 3 1 2 0 1 3 3
3 3 1 3
6 3 0 2 3 0 2
32 3 3 1 3 0 3 0 1 3 0 2 1 3 1 3 3 3 1 3 3 1 2 1 1 3 0 1 3 3 3 1 3
4 3 1 1 1
1 3
2 3 3
2 3 3
14 3 3 1 3 3 3 1 3 0 3 0 1 3 3
11 3 1 1 2 3 0 1 2 0 2 3
3 3 3 0
18 3 0 3 1 3 0 3 1 3 0 2 3 0 0 1 1 1 3
9 3 1 3 0 3 3 3 0 3
6 3 1 3 0 1 3
3 3 3 2
3 3 3 0
7 3 3 0 1 2 3 0
6 3 0 3 1 3 3
6 3 3 0 0 1 3
2 3 3
2 3 3
23 3 2 0 3 0 2 0 2 3 0 2 0 1 3 3 0 3 0 1 3 3 0 1
18 3 1 1 3 1 2 0 2 0 3 0 1 3 3 0 3 0 1
26 3 0 3 0 0 1 3 3 1 3 3 1 0 0 1 3 3 1 3 0 1 2 0 3 0 2
2 3 3
2 3 3
10 3 0 1 3 3 3 2 0 0 0
3 3 3 0
18 3 3 1 3 3 3 1 3 3 1 3 3 0 2 1 1 3 0
3 3 3 2
12 3 3 2 3 1 2 0 1 2 0 3 3
11 3 1 3 0 0 0 0 1 2 0 3
14 3 1 3 0 2 0 1 2 1 0 3 2 1 3
2 3 3
2 3 3
10 3 0 3 0 0 2 0 1 3 1
6 3 0 3 1 2 3
2 3 3
6 3 1 1 3 0 3
10 3 0 3 3 0 2 2 0 3 0
3 3 1 3
5 3 3 0 2 3
1 3
8 3 0 3 3 1 3 3 3
6 3 3 2 3 1 0
9 3 3 0 0 3 3 0 3 1
6 3 1 1 3 3 3
1 3
20 3 0 3 0 3 0 1 1 3 3 3 1 3 0 3 0 1 3 3 3
8 3 3 1 1 3 0 3 0
3 3 3 0
1 3
7 3 1 3 0 2 0 3
2 3 3
3 3 0 3
11 3 0 3 1 2 1 1 1 2 1 3
7 3 0 3 3 0 2 1
12 3 3 0 2 0 1 3 3 0 1 2 3
2 3 3
7 3 3 3 1 1 1 3
10 3 0 3 3 3 0 3 3 0 3
1 3
7 3 0 3 1 2 0 3
2 3 3
6 3 0 3 3 3 0
3 3 1 3
4 3 3 0 0
10 3 3 0 2 0 3 0 3 3 2
9 3 0 0 1 2 3 1 3 3
2 3 3
9 3 3 1 3 3 1 3 0 0
25 3 3 0 1 1 1 1 1 2 0 3 0 3 0 3 3 0 2 0 3 1 2 2 0 3
8 3 3 2 3 1 1 1 1
21 3 1 1 0 0 1 3 3 3 0 1 3 3 0 1 3 3 1 3 0 2
11 3 3 0 2 0 3 0 1 0 0 1
3 3 3 2
6 3 0 3 1 3 3
2 3 0
9 3 3 0 1 2 0 3 0 3
10 3 3 1 3 3 0 2 1 3 1
7 3 3 1 0 3 1 1
3 3 1 3
9 3 0 3 0 1 1 3 1 3
10 3 1 1 3 0 1 1 1 1 1
5 3 3 1 3 3
24 3 1 1 3 1 3 0 0 0 2 0 3 0 0 3 0 0 2 0 3 1 1 3 0
6 3 3 1 3 3 3
6 3 0 3 0 2 3
2 3 3
16 3 3 1 3 0 1 3 3 0 1 2 2 0 3 1 1
3 3 1 1
4 3 0 3 0
1 3
3 3 3 0
3 3 0 1
6 3 2 0 3 0 0
3 3 3 0
2 3 3
5 3 3 2 3 0
12 3 3 0 0 3 3 0 1 3 0 2 3
8 3 0 1 2 2 0 3 0
6 3 1 1 3 0 0
2 3 3
22 3 3 0 2 2 0 3 0 0 0 0 0 0 3 0 1 3 3 1 2 1 1
2 3 3
22 3 0 2 3 0 0 1 3 1 1 3 3 3 3 3 3 0 3 0 2 0 3
4 3 2 0 3
8 3 0 3 0 1 3 1 0
3 3 0 3
3 3 3 0
3 3 3 0
3 3 1 3
10 3 0 2 3 2 0 1 2 3 0
5 3 3 1 3 3
21 3 0 3 0 2 3 0 0 1 3 0 1 1 3 1 1 0 2 2 0 0
2 3 3
4 3 0 1 1
4 3 3 2 1
3 3 1 3
2 3 3
3 3 0 1
7 3 0 3 0 0 3 3
8 3 3 0 1 3 3 3 0
8 3 1 1 1 1 1 3 0
4 3 3 1 3
2 3 3
22 3 0 3 1 2 1 0 2 0 2 3 0 2 0 3 0 2 2 2 1 3 0
17 3 3 0 2 2 3 0 1 2 3 1 2 3 0 3 0 3
3 3 0 1
11 3 1 1 3 3 3 2 0 1 3 2
6 3 3 2 0 1 0
10 3 3 0 0 0 3 3 3 0 3
6 3 1 1 3 3 3
3 3 0 3
5 3 0 2 1 3
4 3 3 1 3
9 3 1 1 1 1 3 1 3 0
18 3 0 3 0 3 1 2 2 0 2 0 2 3 0 3 0 2 3
23 3 1 3 0 2 3 1 3 3 3 0 2 1 2 1 3 3 0 0 3 0 0 3
5 3 0 3 0 2
5 3 2 0 1 3
6 3 0 0 0 2 1
1 3
6 3 1 3 0 2 1
3 3 3 2
4 3 3 1 0
4 3 0 2 3
9 3 0 2 1 3 0 2 0 3
2 3 3
8 3 0 3 3 3 1 1 3
2 3 3
2 3 3
9 3 3 2 1 3 2 2 0 3
9 3 1 3 0 1 1 2 1 3
14 3 3 0 1 1 0 1 3 0 1 2 2 0 3
7 3 0 2 1 3 0 0
17 3 3 1 0 1 3 3 0 1 3 3 0 3 3 3 0 3
3 3 0 3
6 3 0 3 1 0 3
1 3
4 3 0 3 0
4 3 0 2 3
15 3 0 3 0 3 0 2 3 0 2 3 1 3 3 0
2 3 3
6 3 1 1 3 0 2
2 3 0
6 3 0 3 3 0 0
4 3 3 1 0
2 3 3
7 3 2 2 3 1 1 3
14 3 3 1 3 3 0 3 1 3 0 3 0 3 2
12 3 0 3 0 1 3 3 1 3 0 3 3
3 3 1 3
2 3 3
3 3 1 3
10 3 0 3 1 2 3 0 1 0 1
4 3 1 0 3
20 3 0 3 1 2 1 2 0 3 0 1 2 1 0 0 3 1 2 1 0
2 3 3
4 3 1 3 0
5 3 3 3 0 3
13 3 0 3 0 1 3 3 0 3 0 3 1 2
3 3 0 3
10 3 3 0 1 1 2 0 3 3 2
1 3
7 3 3 1 0 3 3 2
3 3 0 3
2 3 0
3 3 3 2
7 3 0 1 2 2 0 3
6 3 0 2 1 1 3
15 3 0 2 1 1 3 0 2 3 2 1 2 0 2 0
3 3 0 3
11 3 1 1 3 3 1 3 0 0 0 1
2 3 3
3 3 1 3
2 3 3
8 3 1 3 1 3 3 1 2
3 3 3 3
4 3 3 2 3
1 3
2 3 3
18 3 1 3 0 1 0 0 1 3 3 1 1 3 3 0 0 1 3
10 3 0 3 1 2 3 0 0 0 1
9 3 0 3 1 2 2 0 2 3
1 3
16 3 0 2 1 3 1 3 3 1 3 0 3 0 1 3 3
14 3 0 3 3 1 3 3 1 3 3 0 0 1 3
9 3 0 3 0 1 1 1 1 0
4 3 0 3 0
2 3 3
2 3 0
29 3 3 0 0 0 3 3 3 0 1 0 3 2 0 3 0 1 3 0 3 3 3 1 0 1 3 3 0 3
4 3 1 1 3
4 3 0 3 0
7 3 1 0 1 1 3 0
7 3 1 3 1 2 3 3
11 3 3 1 3 3 3 0 1 1 1 1
2 3 3
8 3 1 3 0 0 0 1 1
11 3 0 3 1 2 1 2 0 3 3 0
3 3 1 3
1 3
12 3 3 1 3 3 3 0 2 0 3 0 2
6 3 3 1 3 3 3
22 3 3 0 0 3 3 2 1 1 3 0 3 0 1 1 3 3 0 3 0 2 3
1 3
3 3 0 3
6 3 3 2 0 2 1
3 3 3 0
15 3 3 0 1 1 0 1 2 3 0 2 1 1 2 0
5 3 0 3 3 0
33 3 1 3 1 3 3 1 2 1 3 3 3 3 3 1 2 1 1 1 3 0 3 1 2 0 0 1 3 1 2 3 3 1
8 3 0 3 3 0 0 0 2
13 3 0 0 2 3 0 2 0 2 2 3 0 3
2 3 0
5 3 1 3 1 3
29 3 0 3 1 0 1 3 1 2 1 1 2 3 0 3 3 0 2 2 0 3 1 2 2 0 3 3 0 0
10 3 3 1 3 3 1 3 0 3 3
17 3 1 3 0 2 0 2 3 1 1 3 3 0 0 0 1 1
10 3 0 3 0 1 0 1 2 1 3
13 3 0 3 1 3 0 3 3 0 0 0 1 0
24 3 0 0 3 2 3 1 1 3 1 1 1 2 3 1 3 3 3 0 2 0 3 1 0
8 3 0 3 1 2 1 0 3
15 3 1 3 0 2 1 1 1 3 3 3 0 1 2 0
3 3 0 3
19 3 0 3 3 1 3 3 3 0 1 3 3 3 3 2 0 2 2 0
3 3 1 3
13 3 1 1 3 3 3 1 2 3 1 3 0 0
1 3
6 3 0 3 1 3 0
2 3 3
3 3 3 0
5 3 0 3 1 3
7 3 3 3 1 3 0 3
4 3 3 0 2
7 3 1 1 1 1 1 1
3 3 3 0
4 3 0 3 3
2 3 3
3 3 0 3
5 3 1 1 3 0
3 3 1 3
4 3 3 0 0
3 3 1 1
2 3 3
15 3 3 0 1 2 1 3 1 3 3 2 1 1 0 1
4 3 3 0 1
4 3 1 1 3
9 3 0 3 0 0 3 0 1 2
6 3 3 2 0 0 2
1 3
5 3 0 1 3 3
7 3 3 0 2 1 2 0
3 3 1 3
8 3 0 3 3 0 1 2 3
10 3 0 3 0 2 0 0 0 1 3
3 3 3 0
16 3 1 1 3 0 2 1 1 1 1 1 1 3 1 3 0
3 3 1 3
7 3 0 3 0 3 0 1
1 3
2 3 3
2 3 3
4 3 0 3 3
1 3
28 3 1 3 0 2 2 0 1 1 3 1 3 3 3 0 0 1 3 0 0 0 1 1 0 2 0 3 0
5 3 1 1 3 3
22 3 0 3 1 2 2 0 0 0 1 3 3 0 0 3 0 1 3 3 0 3 3
5 3 1 2 3 3
4 3 0 3 3
10 3 3 1 3 3 1 0 2 0 3
10 3 3 0 1 0 1 3 3 3 0
2 3 3
9 3 0 3 1 2 2 0 1 1
1 3
8 3 3 1 2 1 3 0 0
3 3 3 2
10 3 0 3 0 1 1 1 3 2 3
5 3 1 1 1 2
5 3 1 3 3 3
3 3 0 3
3 3 3 2
4 3 1 3 0
3 3 3 2
6 3 1 1 3 3 3
3 3 3 0
1 3
6 3 3 1 3 3 3
14 3 0 3 0 1 3 3 3 0 2 0 3 0 1
3 3 3 2
4 3 0 3 0
7 3 1 3 0 1 1 0
4 3 0 2 3
2 3 0
5 3 2 0 3 0
29 3 3 2 0 2 3 2 2 0 0 3 0 2 0 3 0 2 3 0 2 1 1 1 1 1 1 1 1 3
11 3 0 1 2 0 3 0 1 2 0 3
4 3 3 0 2
5 3 1 1 3 0
8 3 3 1 3 3 3 1 2
4 3 2 0 3
31 3 0 3 0 3 0 2 3 0 1 1 2 3 0 1 0 1 3 3 0 3 0 1 0 3 3 1 2 1 1 0
2 3 3
34 3 0 3 2 0 1 3 1 3 3 0 3 0 1 0 3 3 0 3 3 1 0 1 0 0 1 3 3 3 1 3 3 1 3
2 3 3
3 3 3 0
3 3 0 3
4 3 3 0 0
14 3 3 0 1 1 2 0 3 1 3 0 3 0 3
2 3 3
9 3 1 1 1 1 1 3 3 3
3 3 0 1
5 3 1 3 1 3
5 3 0 3 1 3
6 3 1 0 3 3 3
3 3 0 3
1 3
6 3 0 3 0 3 3
3 3 3 2
12 3 0 3 3 1 3 3 3 0 2 0 3
3 3 1 3
5 3 0 3 0 3
11 3 0 3 0 2 3 1 1 1 2 0
2 3 3
7 3 0 3 0 2 1 3
4 3 0 2 3
22 3 1 1 3 3 0 1 0 0 1 2 3 0 0 1 3 0 1 0 3 3 2
7 3 1 1 3 1 3 0
1 3
1 3
7 3 3 2 3 0 0 3
2 3 3
8 3 0 3 3 0 2 0 3
8 3 3 0 1 2 3 2 0
6 3 3 1 1 0 3
5 3 1 3 1 0
4 3 1 3 0
2 3 0
13 3 0 1 3 3 3 1 3 3 1 2 0 3
4 3 3 2 0
2 3 3
7 3 2 0 3 0 1 1
4 3 2 0 3
7 3 3 1 1 1 3 0
3 3 0 3
4 3 0 3 3
4 3 3 2 3
9 3 0 3 1 3 0 1 1 0
4 3 1 1 3
5 3 1 0 3 3
1 3
10 3 0 2 3 0 2 1 2 0 1
7 3 0 3 1 3 0 2
22 3 0 3 0 1 1 3 0 2 1 2 0 3 0 3 0 2 0 1 1 1 3
6 3 1 3 2 1 3
4 3 0 2 3
16 3 3 1 3 3 1 3 3 0 3 1 2 1 1 1 0
13 3 3 2 0 2 3 3 1 3 0 0 2 3
9 3 0 3 1 3 3 0 1 3
17 3 3 1 3 3 0 1 3 3 1 2 1 1 3 1 0 2
2 3 3
2 3 3
2 3 3
10 3 3 2 0 0 3 3 1 1 1
12 3 3 1 2 1 1 1 1 1 2 0 3
3 3 2 2
1 3
3 3 3 1
16 3 1 1 3 1 3 1 3 0 1 3 3 1 2 0 3
3 3 0 3
3 3 3 0
4 3 3 0 0
7 3 1 2 0 1 0 1
15 3 0 1 3 2 2 3 0 1 2 0 1 0 3 3
7 3 1 3 0 2 3 1
9 3 0 3 0 1 3 3 1 3
23 3 0 3 1 2 1 1 2 0 3 1 0 1 3 3 0 3 3 0 1 3 2 3
5 3 3 0 2 0
15 3 0 3 1 0 1 3 2 3 1 3 3 2 1 0
3 3 1 3
3 3 1 3
5 3 0 3 1 3
6 3 0 3 0 2 2
4 3 1 3 0
4 3 1 3 0
8 3 0 3 1 2 1 1 3
4 3 1 1 3
11 3 2 0 3 0 1 1 2 0 3 3
2 3 3
2 3 0
2 3 3
3 3 0 3
5 3 3 0 0 0
3 3 1 3
20 3 0 3 1 3 0 3 0 1 3 3 1 2 3 0 0 1 3 0 0
5 3 1 1 1 3
3 3 3 2
27 3 1 0 3 3 0 1 2 1 1 1 1 1 1 1 1 2 0 3 0 1 3 3 0 3 0 2
8 3 0 1 2 0 1 3 0
2 3 3
5 3 3 1 2 3
10 3 3 1 3 3 1 2 1 1 0
7 3 0 1 3 3 3 1
1 3
6 3 3 0 1 2 3
20 3 3 1 3 3 1 0 1 3 3 0 1 3 3 0 1 1 0 2 3
5 3 1 1 3 0
12 3 0 3 0 3 0 1 2 0 1 3 0
8 3 0 3 0 2 0 3 0
5 3 3 1 0 3
4 3 3 1 3
21 3 0 3 3 2 0 2 2 2 3 1 2 2 3 1 3 2 0 1 3 0
9 3 1 1 1 1 3 3 0 0
37 3 3 1 3 3 3 0 2 0 3 0 1 3 3 0 3 3 2 3 0 3 1 2 2 0 3 0 3 0 1 3 3 0 3 3 2 1
4 3 1 3 0
11 3 0 2 3 0 1 1 1 2 0 3
2 3 3
10 3 0 3 1 0 1 0 1 0 2
16 3 0 3 3 1 0 0 3 3 0 3 0 2 1 3 2
3 3 0 3
6 3 0 3 0 2 1
4 3 3 1 2
14 3 0 3 0 3 0 3 1 2 1 1 0 3 3
7 3 0 2 1 1 3 0
14 3 1 0 0 0 1 3 3 0 1 1 3 3 2
12 3 0 3 0 1 3 3 1 0 1 0 0
2 3 0
5 3 0 3 0 3
6 3 0 3 1 0 2
2 3 3
5 3 1 3 1 3
10 3 3 1 3 3 1 2 2 0 3
7 3 3 1 3 3 0 2
3 3 1 3
7 3 3 1 3 3 3 3
5 3 1 0 3 1
9 3 1 1 1 1 1 1 1 3
6 3 2 0 1 3 0
2 3 3
2 3 3
10 3 3 0 1 3 0 1 2 3 3
2 3 0
10 3 1 1 3 1 3 1 0 1 3
6 3 1 1 3 1 3
4 3 1 3 0
11 3 3 0 2 0 3 1 2 1 1 3
1 3
12 3 3 1 2 3 0 3 1 3 3 0 2
4 3 1 3 0
9 3 1 3 0 2 1 2 0 1
8 3 3 1 3 0 3 3 0
2 3 1
4 3 0 3 3
7 3 0 3 0 1 2 3
11 3 0 2 3 3 3 3 0 1 0 3
2 3 3
3 3 0 3
4 3 0 3 0
3 3 0 1
5 3 3 0 1 0
2 3 3
1 3
15 3 1 3 0 0 3 3 1 0 1 3 3 1 2 3
1 3
1 3
8 3 0 3 0 2 0 3 0
4 3 3 2 0
3 3 0 3
1 3
20 3 0 3 1 3 0 3 0 1 2 2 0 3 2 0 1 3 1 3 3
6 3 0 3 1 0 2
3 3 1 3
3 3 1 3
8 3 0 3 1 3 2 0 3
2 3 3
6 3 3 0 2 0 3
2 3 3
6 3 3 0 1 0 2
4 3 3 0 2
6 3 3 1 3 1 2
9 3 3 1 0 2 3 1 1 2
1 3
21 3 0 3 0 1 3 3 1 2 2 3 1 3 3 0 3 0 0 2 1 0
3 3 0 3
25 3 0 2 3 1 3 3 0 3 1 0 1 2 1 1 1 2 3 1 3 3 0 1 2 3
3 3 3 0
3 3 0 3
10 3 0 3 0 1 1 3 2 1 0
8 3 3 1 3 3 0 2 3
6 3 1 1 1 1 3
7 3 0 3 0 1 3 3
3 3 1 0
16 3 0 3 3 3 3 0 3 3 3 2 3 1 2 0 1
6 3 0 3 1 2 3
13 3 0 3 1 3 0 2 1 1 3 1 3 0
2 3 3
7 3 3 1 1 1 1 3
7 3 3 0 1 1 1 3
16 3 3 1 1 1 3 1 1 1 1 3 0 0 3 0 0
6 3 1 3 0 2 1
3 3 3 0
3 3 3 0
3 3 0 3
15 3 1 3 1 3 3 3 1 2 1 3 1 1 0 0
11 3 3 0 1 1 1 1 2 0 2 3
2 3 3
2 3 0
2 3 3
7 3 1 3 0 0 1 3
11 3 0 3 1 3 0 2 3 0 0 0
6 3 3 0 2 3 3
3 3 3 2
7 3 3 0 2 0 3 0
5 3 0 3 0 2
8 3 0 3 0 1 2 3 0
4 3 3 0 0
2 3 1
2 3 0
2 3 3
3 3 1 3
3 3 1 3
17 3 3 1 3 3 2 0 0 3 0 2 3 2 3 1 2 3
24 3 0 2 3 0 1 2 0 3 0 2 1 0 1 3 3 1 2 1 0 1 3 0 0
3 3 3 0
2 3 1
8 3 0 3 1 2 0 3 0
5 3 3 0 1 0
3 3 3 0
10 3 0 3 3 0 2 2 0 1 3
3 3 0 2
5 3 1 1 1 1
3 3 3 0
32 3 0 3 0 1 3 3 3 0 2 0 2 3 0 2 1 3 3 3 0 1 1 3 0 2 1 1 1 3 3 0 2
3 3 3 2
3 3 1 3
8 3 0 3 1 3 3 0 0
4 3 0 3 0
9 3 3 1 3 3 1 2 0 3
14 3 0 3 1 2 2 0 3 0 3 1 0 1 0
17 3 3 1 3 3 0 2 1 3 0 2 0 1 2 0 1 2
4 3 0 3 3
13 3 3 0 0 0 1 3 3 3 0 1 3 3
14 3 3 2 1 3 3 0 3 3 0 0 1 3 0
13 3 1 1 1 1 1 1 3 0 0 1 1 3
6 3 3 0 0 1 3
5 3 1 1 3 3
5 3 1 3 0 0
9 3 1 0 3 3 2 0 1 3
2 3 1
8 3 1 3 1 1 1 3 0
22 3 3 1 3 3 1 1 0 1 0 3 3 0 1 1 3 3 2 2 0 3 3
1 3
3 3 3 2
12 3 3 1 3 3 0 2 1 3 0 1 3
5 3 1 0 3 3
3 3 3 2
3 3 0 3
4 3 1 1 3
26 3 0 3 3 0 1 1 1 1 3 2 1 2 3 1 3 0 3 1 2 3 1 3 3 0 3
2 3 3
25 3 3 0 2 3 0 3 0 2 3 0 1 1 3 2 1 3 2 3 1 3 3 0 2 3
13 3 1 3 1 1 3 0 3 3 3 3 1 0
21 3 0 3 0 3 0 1 2 1 2 0 3 0 1 3 3 0 3 1 1 3
3 3 1 3
3 3 0 2
4 3 1 3 0
10 3 3 1 3 1 3 3 0 2 3
8 3 0 3 1 0 2 1 0
4 3 0 3 3
3 3 3 1
6 3 1 3 0 0 3
5 3 0 3 1 3
2 3 3
2 3 3
5 3 0 3 0 2
12 3 0 3 0 2 3 1 1 3 3 3 1
8 3 0 3 1 2 1 1 1
24 3 1 1 1 3 0 1 3 3 3 0 3 0 1 2 3 0 3 1 0 1 3 3 0
5 3 0 2 3 0
3 3 3 0
12 3 0 2 3 1 0 2 1 1 1 1 3
5 3 3 0 0 0
2 3 0
25 3 1 3 0 2 2 0 3 1 0 1 3 1 3 0 1 2 0 3 1 0 1 3 3 0
18 3 1 3 2 0 2 3 1 0 1 3 3 1 3 0 0 1 3
14 3 0 3 1 2 1 2 0 3 0 1 0 1 3
2 3 3
3 3 0 3
2 3 3
6 3 0 3 1 0 2
2 3 3
19 3 3 1 2 1 0 0 1 1 3 3 0 2 0 3 1 2 0 3
1 3
14 3 0 2 3 0 1 1 1 2 0 3 0 0 3
9 3 1 1 3 0 0 1 3 0
18 3 0 2 0 0 0 3 3 3 3 3 1 3 1 3 0 0 0
9 3 1 1 3 1 3 0 2 3
4 3 0 2 3
2 3 3
9 3 1 1 1 1 3 1 3 3
2 3 3
18 3 3 1 0 2 3 0 3 1 3 1 1 3 1 1 0 0 3
4 3 0 1 0
3 3 1 2
2 3 3
4 3 0 3 3
11 3 0 2 3 3 0 3 0 1 0 2
1 3
2 3 0
10 3 0 3 1 2 0 3 0 1 1
5 3 0 3 1 2
8 3 3 0 3 0 3 1 3
5 3 3 1 3 3
1 3
7 3 0 3 1 2 0 3
12 3 3 1 3 3 3 0 1 3 3 0 3
17 3 0 3 1 2 1 3 0 2 3 1 3 3 3 1 1 3
5 3 0 3 0 1
1 3
21 3 3 1 3 3 0 3 0 1 3 3 1 2 3 0 1 2 3 2 0 0
52 3 0 3 1 0 1 0 1 3 3 0 2 0 3 1 3 3 0 1 3 3 0 3 0 1 3 3 0 3 3 1 3 3 3 1 1 1 1 1 2 1 3 0 1 1 1 1 2 0 3 3 3
6 3 0 1 3 3 3
6 3 0 3 0 2 3
4 3 3 0 1
3 3 1 3
3 3 3 0
17 3 3 0 1 1 3 2 1 1 2 3 1 3 0 3 0 2
6 3 0 2 3 0 3
5 3 3 1 1 3
11 3 3 0 1 2 3 1 3 3 0 3
7 3 1 2 0 2 1 3
9 3 0 3 1 0 1 3 3 0
4 3 0 3 0
3 3 1 1
5 3 3 0 2 1
3 3 1 0
18 3 0 3 0 0 3 1 1 1 0 2 2 3 0 1 3 3 3
4 3 0 3 0
8 3 0 3 1 3 1 3 2
5 3 0 2 1 3
3 3 0 3
9 3 0 3 1 0 2 1 2 3
6 3 0 3 1 2 3
4 3 3 0 0
14 3 0 3 1 0 1 2 1 3 3 1 0 3 3
4 3 3 0 2
7 3 0 3 1 2 1 3
15 3 0 3 0 2 1 1 0 2 0 2 0 3 1 3
6 3 1 3 0 0 0
9 3 0 2 0 1 3 3 0 3
12 3 3 1 0 2 1 3 3 3 0 1 0
24 3 3 1 3 0 1 2 1 1 1 1 1 1 1 1 3 1 1 0 1 3 3 3 0
6 3 3 2 0 2 3
15 3 0 3 3 1 3 0 1 3 3 1 0 1 2 3
4 3 1 0 0
8 3 1 1 1 3 1 3 3
1 3
12 3 3 1 3 3 1 2 3 0 0 1 3
29 3 0 3 1 2 1 1 3 3 1 3 2 3 1 2 2 3 0 2 2 3 0 2 3 1 3 3 1 2
2 3 3
5 3 0 3 0 2
2 3 3
6 3 0 3 1 3 3
10 3 3 0 1 1 2 0 3 0 3
4 3 0 3 2
2 3 3
4 3 1 3 0
9 3 0 3 0 1 3 3 1 2
3 3 0 1
2 3 3
14 3 0 3 0 2 3 0 2 3 1 2 1 3 3
28 3 0 0 2 3 1 3 3 1 0 2 3 1 3 0 0 3 0 1 1 1 1 1 1 1 3 1 3
4 3 1 3 0
6 3 3 0 2 3 3
2 3 3
3 3 3 3
5 3 0 3 0 3
26 3 3 0 3 3 0 1 2 1 1 0 2 0 1 3 3 1 3 0 3 1 3 3 3 0 1
3 3 0 3
2 3 3
8 3 0 1 2 1 3 2 0
3 3 1 3
3 3 0 3
5 3 3 1 3 3
9 3 3 0 1 2 0 3 1 3
11 3 3 2 0 1 2 1 3 0 2 3
11 3 0 3 1 2 2 0 3 3 0 2
1 3
2 3 3
3 3 1 3
14 3 0 3 3 1 3 3 1 2 0 3 0 0 3
2 3 0
3 3 3 0
3 3 0 1
3 3 0 3
4 3 0 3 3
5 3 0 2 2 3
3 3 0 1
3 3 0 1
11 3 0 1 3 3 3 0 2 0 2 3
2 3 2
6 3 3 0 1 1 1
5 3 1 3 0 0
3 3 1 3
1 3
21 3 0 3 1 2 0 1 3 1 3 1 1 1 2 0 3 3 1 2 2 3
1 3
4 3 3 0 0
3 3 3 0
16 3 0 2 1 0 2 0 0 0 1 1 3 0 2 1 2
6 3 0 0 2 1 3
13 3 3 0 1 1 0 1 3 1 2 3 0 0
22 3 1 3 1 3 3 1 3 0 1 0 1 3 2 3 0 3 0 1 3 3 0
15 3 0 3 0 0 3 0 1 2 0 2 0 2 3 0
10 3 0 2 3 0 2 3 2 1 2
4 3 0 3 3
4 3 0 3 3
4 3 3 0 2
1 3
6 3 1 1 1 1 3
4 3 3 2 3
1 3
2 3 3
3 3 0 3
14 3 0 3 0 3 3 3 1 3 3 1 2 0 0
4 3 0 3 1
8 3 3 0 0 3 3 3 3
2 3 0
4 3 3 0 2
9 3 3 2 3 2 0 3 0 0
2 3 3
8 3 1 3 1 1 2 1 0
3 3 3 0
2 3 3
11 3 0 3 0 1 3 3 3 0 1 1
14 3 0 3 0 1 3 2 0 1 2 1 3 0 2
10 3 0 3 1 0 1 0 1 3 3
4 3 3 0 2
3 3 1 3
11 3 0 3 1 3 0 1 3 3 0 3
1 3
2 3 3
3 3 0 1
19 3 2 0 3 1 3 3 3 1 3 3 0 3 0 3 0 0 0 2
12 3 3 0 0 0 1 0 1 2 1 3 3
7 3 3 0 1 1 1 3
3 3 0 1
8 3 0 3 1 3 0 3 3
25 3 0 3 1 0 1 3 3 1 3 0 3 0 1 2 1 2 0 3 0 1 2 3 1 2
3 3 1 3
4 3 3 0 0
8 3 0 2 3 1 0 1 3
25 3 0 3 3 0 3 3 1 3 0 3 1 2 1 1 1 1 2 0 2 3 1 0 0 0
1 3
3 3 0 3
10 3 0 1 0 1 3 3 1 3 0
2 3 3
9 3 3 1 1 1 1 3 1 3
12 3 3 1 3 3 1 2 0 3 0 0 3
5 3 1 1 3 0
5 3 0 3 1 3
4 3 0 2 3
2 3 3
42 3 0 1 2 1 2 1 3 3 3 1 3 3 3 0 1 0 1 3 3 3 0 3 3 0 1 3 2 1 1 1 2 0 3 3 0 0 1 3 0 0 3
8 3 0 3 1 0 1 3 3
4 3 3 0 0
9 3 0 3 3 0 1 2 3 0
21 3 0 3 1 2 2 0 3 3 0 1 1 2 0 3 3 1 1 1 3 0
13 3 1 1 3 1 1 1 1 1 1 1 1 1
4 3 1 3 0
8 3 0 3 1 3 1 0 2
2 3 3
2 3 3
5 3 1 3 0 2
6 3 1 2 1 3 3
6 3 0 3 0 3 0
2 3 3
2 3 3
8 3 0 1 3 3 2 0 3
2 3 1
5 3 1 1 1 3
11 3 0 3 0 3 1 0 1 3 3 3
7 3 3 1 2 1 2 0
3 3 3 0
3 3 1 3
27 3 0 3 1 2 1 1 1 2 3 1 3 3 3 3 0 1 1 2 3 1 3 3 0 0 1 2
9 3 2 0 3 0 2 1 1 3
6 3 2 0 3 0 2
3 3 0 1
8 3 3 0 2 0 0 2 3
12 3 3 3 1 2 1 1 2 0 2 3 0
4 3 0 3 0
4 3 0 3 1
8 3 3 1 0 1 0 1 0
13 3 0 2 2 1 1 1 1 1 0 1 1 2
2 3 3
6 3 0 1 3 3 3
5 3 0 3 1 3
5 3 1 3 0 2
4 3 2 0 3
11 3 3 0 1 2 1 3 0 0 1 3
3 3 3 0
2 3 3
16 3 0 3 1 3 0 2 3 1 3 1 3 0 0 1 3
2 3 3
2 3 3
1 3
10 3 0 3 0 1 3 3 1 3 1
5 3 0 2 3 0
9 3 3 1 3 3 1 2 0 3
10 3 3 0 1 2 1 1 2 0 2
12 3 0 3 1 2 3 1 3 3 0 0 2
5 3 3 0 0 0
4 3 1 3 0
5 3 0 3 3 0
11 3 3 1 3 3 3 0 1 1 2 0
3 3 0 3
5 3 3 1 3 3
25 3 0 3 0 3 0 3 0 1 3 2 3 3 3 3 3 1 3 3 0 3 1 2 0 3
22 3 0 3 1 3 3 0 2 1 3 0 2 0 1 3 3 1 2 1 1 1 0
2 3 3
9 3 3 0 2 0 1 0 0 1
3 3 0 3
6 3 3 0 1 2 3
4 3 1 3 0
2 3 0
3 3 3 1
4 3 0 3 0
2 3 3
2 3 3
2 3 3
7 3 1 2 1 1 3 3
10 3 3 0 2 2 0 0 3 0 0
8 3 0 3 1 3 1 1 3
5 3 1 1 1 3
27 3 0 3 0 1 3 3 3 3 0 3 1 2 1 2 3 1 3 3 0 3 0 1 3 3 1 0
5 3 1 3 0 2
7 3 3 3 0 1 1 0
7 3 1 1 3 1 3 0
3 3 1 2
16 3 0 3 0 2 0 0 2 0 3 1 2 2 0 3 0
2 3 3
7 3 1 3 3 1 3 3
8 3 0 3 1 2 2 0 3
6 3 3 0 3 3 0
4 3 1 3 0
14 3 3 0 1 1 1 1 1 1 2 0 2 2 3
10 3 0 3 3 3 0 2 1 2 0
2 3 3
2 3 3
3 3 1 3
2 3 3
7 3 3 2 0 2 3 0
2 3 3
4 3 3 0 2
15 3 0 2 1 1 2 1 0 1 3 3 3 0 0 1
2 3 3
12 3 3 1 2 3 1 3 3 3 0 2 1
19 3 0 2 3 0 2 3 0 0 1 2 3 0 0 3 2 3 0 3
4 3 2 1 0
5 3 3 1 3 3
13 3 3 1 1 0 1 3 3 3 2 3 0 3
3 3 0 3
5 3 3 0 2 3
3 3 3 1
4 3 3 1 3
6 3 1 1 1 1 3
3 3 0 3
1 3
3 3 0 3
3 3 0 3
6 3 0 3 1 3 3
19 3 0 3 0 3 0 1 3 3 0 1 1 1 3 3 0 0 0 0
2 3 3
7 3 3 2 0 0 1 3
8 3 3 0 2 1 1 0 3
5 3 0 3 3 2
13 3 3 0 2 0 3 1 2 1 1 3 2 1
6 3 1 3 1 3 3
3 3 0 3
2 3 3
3 3 0 3
6 3 0 1 3 3 3
14 3 0 3 0 1 2 0 3 0 0 1 1 3 0
11 3 0 3 1 3 0 1 3 3 1 0
24 3 3 1 2 1 2 0 3 0 1 2 1 1 2 0 3 0 3 0 0 1 2 0 3
8 3 0 2 0 1 0 1 0
7 3 0 0 2 2 0 3
2 3 3
14 3 1 0 3 1 2 0 3 0 1 1 1 3 0
9 3 1 3 0 0 0 3 3 3
10 3 0 1 2 1 2 3 3 0 0
5 3 1 2 0 1
14 3 1 3 0 2 3 1 3 3 3 1 3 3 0
13 3 0 3 0 3 1 2 1 2 0 3 0 2
2 3 3
5 3 1 1 1 3
2 3 3
2 3 3
7 3 0 3 1 2 3 0
2 3 3
5 3 3 1 3 0
4 3 0 3 0
8 3 3 0 2 2 3 1 3
11 3 0 3 0 2 3 0 2 3 1 0
17 3 0 3 0 2 1 0 1 0 3 1 2 3 0 1 1 3
6 3 1 3 0 0 0
4 3 1 3 0
9 3 0 3 1 2 2 3 0 0
2 3 3
10 3 0 3 1 2 0 3 0 0 0
3 3 0 1
22 3 0 3 0 1 2 1 0 1 3 0 1 3 3 0 2 1 3 0 0 3 0
17 3 0 3 1 3 3 2 3 0 1 3 2 1 3 2 1 0
3 3 0 2
2 3 3
1 3
3 3 3 0
3 3 0 3
7 3 1 0 3 3 3 1
10 3 3 1 0 1 0 1 3 0 3
7 3 3 1 2 0 3 3
13 3 1 2 0 0 1 3 0 2 0 3 0 3
17 3 1 3 0 0 0 3 3 3 0 1 0 1 0 1 2 1
8 3 0 2 3 0 0 1 3
6 3 0 3 0 2 3
15 3 3 0 2 0 3 0 1 3 3 0 1 0 2 0
5 3 3 0 2 3
6 3 3 3 0 0 3
6 3 0 2 3 0 1
4 3 0 1 0
7 3 0 3 0 1 0 3
13 3 3 3 1 3 3 3 1 1 2 1 1 3
2 3 0
27 3 1 1 3 1 3 3 1 3 3 1 3 3 3 2 0 1 2 0 3 1 2 1 1 1 0 3
6 3 3 1 3 3 3
2 3 3
6 3 3 0 2 0 3
4 3 3 3 0
7 3 3 1 3 3 0 1
3 3 3 0
3 3 0 3
6 3 0 3 0 1 1
4 3 3 2 0
2 3 3
8 3 0 3 1 3 0 3 0
21 3 3 2 0 0 1 3 3 3 0 1 0 0 1 3 3 0 2 0 0 1
14 3 0 3 0 1 3 3 0 3 0 3 2 0 3
12 3 1 1 0 3 1 3 0 3 3 3 0
2 3 3
2 3 3
13 3 1 1 1 1 1 3 1 3 3 0 1 2
11 3 3 2 3 1 2 0 2 0 1 0
1 3
13 3 3 1 3 3 0 3 3 0 0 1 3 3
13 3 0 3 0 3 0 2 0 1 2 1 1 0
2 3 3
10 3 2 0 0 3 0 2 3 3 0
13 3 0 3 1 0 1 3 3 1 3 0 1 0
4 3 1 3 0
3 3 0 3
4 3 1 2 0
4 3 1 1 3
7 3 3 1 3 0 3 0
13 3 3 0 2 1 0 3 1 2 1 0 3 3
25 3 3 0 2 0 3 3 0 1 2 0 3 1 3 0 2 3 0 0 0 1 1 2 0 3
14 3 0 1 2 3 3 1 3 3 0 3 0 3 3
17 3 3 1 2 1 1 1 3 2 2 0 3 0 2 0 3 0
3 3 1 3
1 3
6 3 3 0 0 3 3
21 3 1 0 3 3 1 0 1 3 3 0 3 0 3 1 3 0 3 1 2 3
3 3 3 0
20 3 3 0 1 2 3 0 0 1 3 0 1 2 3 1 3 3 1 3 0
20 3 0 2 3 1 1 1 1 3 3 0 0 1 3 3 0 1 3 3 3
1 3
16 3 3 0 2 3 2 2 2 0 0 3 1 3 2 0 3
5 3 0 3 0 3
4 3 0 3 3
4 3 0 3 3
4 3 3 0 3
10 3 3 0 3 0 3 1 2 2 3
13 3 1 1 3 0 1 1 1 1 2 0 2 3
25 3 3 0 2 1 3 2 1 0 2 0 2 3 0 2 1 0 3 3 0 1 2 0 3 1
18 3 3 1 1 3 0 2 0 3 0 2 2 2 3 0 1 1 3
4 3 0 3 3
2 3 3
32 3 3 1 3 3 1 2 2 0 2 3 1 3 3 0 1 0 2 3 0 3 1 0 1 2 3 0 2 1 0 3 1
9 3 0 3 0 1 3 3 0 3
3 3 1 3
8 3 0 2 1 3 0 0 0
3 3 3 0
3 3 1 3
9 3 0 3 1 3 0 1 1 3
13 3 0 3 3 1 3 3 1 2 2 0 3 1
7 3 0 3 1 2 0 3
15 3 0 3 1 2 1 1 2 0 3 1 0 2 0 3
7 3 0 3 0 2 0 3
2 3 3
19 3 0 3 1 2 1 2 0 3 1 2 1 2 0 3 1 0 2 3
4 3 0 3 0
2 3 3
3 3 0 3
2 3 3
3 3 1 3
18 3 1 2 0 1 1 1 1 1 1 2 0 3 1 2 1 1 0
7 3 0 3 0 2 3 0
5 3 3 0 0 3
9 3 0 1 1 0 3 3 0 0
1 3
10 3 0 3 0 1 0 0 0 0 3
2 3 3
3 3 3 0
2 3 3
4 3 1 3 0
9 3 3 1 1 3 2 1 1 3
7 3 3 0 0 1 3 0
8 3 0 3 1 3 0 2 3
10 3 3 1 3 3 0 1 0 2 0
12 3 0 3 1 2 0 3 3 1 3 3 3
3 3 3 2
8 3 3 1 3 3 0 1 3
2 3 1
3 3 1 3
2 3 3
4 3 1 3 1
6 3 0 3 3 3 3
11 3 0 3 1 2 1 1 2 0 3 3
2 3 3
8 3 0 3 0 3 1 3 3
5 3 3 1 0 2
10 3 0 3 0 3 1 3 0 1 2
12 3 3 1 0 3 3 3 3 0 3 1 1
5 3 3 1 3 3
10 3 0 1 1 2 3 0 2 1 2
2 3 3
2 3 3
4 3 1 1 3
6 3 1 3 0 0 0
4 3 1 3 0
13 3 3 3 0 0 1 1 3 1 3 3 3 0
3 3 3 0
7 3 2 0 3 0 2 0
6 3 0 1 1 1 1
25 3 3 1 3 3 0 3 0 3 1 0 1 0 2 3 1 1 2 0 3 3 3 0 2 2
2 3 3
1 3
3 3 3 0
6 3 0 3 1 3 0
6 3 3 0 3 3 3
23 3 1 3 0 2 2 0 0 3 0 0 3 3 3 1 3 3 0 0 3 3 1 3
13 3 0 3 0 3 0 3 0 2 1 0 2 0
7 3 3 1 3 3 1 3
5 3 0 3 1 2
8 3 0 3 1 3 0 2 1
22 3 1 3 0 0 0 1 1 3 0 3 0 2 3 0 3 3 0 1 3 1 0
16 3 0 1 3 3 0 3 3 1 3 0 3 3 3 0 2
4 3 1 1 3
7 3 0 3 2 3 3 3
3 3 0 3
3 3 1 3
2 3 1
2 3 3
12 3 0 3 0 2 0 0 1 2 3 0 0
9 3 1 1 3 1 3 3 0 3
3 3 0 3
7 3 3 0 2 1 2 0
4 3 0 1 2
14 3 0 3 0 1 3 3 0 3 1 2 1 1 1
3 3 0 3
4 3 2 0 3
5 3 0 3 0 2
16 3 0 3 0 2 1 1 3 0 3 0 3 2 1 2 1
4 3 0 2 3
2 3 3
4 3 0 3 0
5 3 0 3 3 0
2 3 3
4 3 0 2 3
4 3 1 1 3
3 3 1 3
9 3 1 3 0 0 3 3 0 3
19 3 1 3 1 3 3 1 3 1 3 3 1 1 0 3 1 3 3 3
1 3
5 3 1 3 2 0
12 3 1 0 3 3 0 2 0 0 1 1 3
16 3 0 3 0 1 0 0 2 3 1 2 1 3 1 2 3
8 3 1 3 0 1 1 1 0
8 3 0 3 3 1 1 3 3
3 3 1 2
11 3 0 1 2 0 3 0 1 3 3 1
2 3 3
3 3 0 3
4 3 2 0 3
5 3 0 3 0 2
24 3 1 3 1 3 3 0 3 0 1 2 3 3 0 0 0 1 0 1 2 3 1 3 0
12 3 0 3 1 0 1 3 3 0 3 0 3
3 3 0 3
1 3
1 3
1 3
9 3 0 3 0 1 2 1 1 0
1 3
17 3 3 3 1 3 0 3 3 1 3 3 3 1 2 1 1 3
5 3 1 1 3 3
7 3 0 3 1 2 3 0
3 3 2 0
1 3
6 3 0 3 1 3 0
3 3 0 3
10 3 0 3 1 0 1 3 3 0 3
8 3 0 3 0 3 1 3 0
11 3 1 3 1 3 3 1 2 1 2 0
7 3 0 2 3 0 0 0
10 3 3 1 2 3 3 1 3 3 3
3 3 0 3
11 3 0 3 0 3 0 3 0 3 0 3
2 3 3
3 3 1 2
3 3 0 3
12 3 0 2 3 1 3 3 3 0 1 0 3
1 3
3 3 0 3
6 3 1 1 1 1 3
5 3 3 0 2 0
8 3 0 3 0 1 3 3 0
16 3 0 3 0 1 3 3 3 0 3 3 0 3 3 0 1
4 3 1 3 2
2 3 3
9 3 0 3 0 2 3 3 3 0
11 3 3 1 3 3 0 3 0 2 0 3
2 3 3
6 3 0 3 0 1 3
5 3 0 1 0 0
12 3 3 1 0 1 3 3 0 1 3 3 3
9 3 3 0 2 0 3 1 3 3
16 3 0 3 0 3 1 3 3 1 3 3 0 1 1 1 1
28 3 3 0 2 3 3 0 2 0 3 1 0 1 1 3 1 1 1 1 1 1 3 3 0 1 3 3 3
6 3 1 1 3 0 0
3 3 0 1
21 3 0 3 1 2 2 0 3 0 2 3 0 0 1 3 0 2 2 0 0 3
11 3 3 1 3 3 1 2 1 3 0 2
7 3 0 3 0 3 3 3
21 3 0 3 0 2 2 3 0 3 0 1 2 1 3 3 3 0 2 2 0 3
8 3 0 3 1 2 2 0 3
6 3 0 3 1 2 3
11 3 3 1 3 3 0 1 3 3 1 3
14 3 0 3 0 0 2 3 0 0 1 1 3 0 2
6 3 3 1 3 3 3
6 3 3 3 2 0 1
17 3 3 0 1 1 3 2 2 0 3 0 1 3 1 3 0 2
6 3 3 0 0 1 3
8 3 0 3 1 2 0 1 3
8 3 3 1 3 3 3 0 3
2 3 1
6 3 1 3 1 3 3
9 3 3 0 2 0 1 1 2 3
11 3 0 2 2 3 0 0 3 0 0 2
2 3 3
13 3 0 3 0 1 3 3 0 3 0 1 2 3
7 3 0 2 3 3 3 3
5 3 1 0 1 3
6 3 0 3 1 3 3
8 3 0 3 1 1 1 1 3
4 3 3 0 2
3 3 3 3
4 3 0 3 1
3 3 0 3
16 3 0 3 0 0 3 0 1 3 3 3 1 2 1 1 0
2 3 3
2 3 3
6 3 0 3 0 1 3
2 3 3
12 3 3 1 3 3 3 0 1 1 2 0 2
2 3 3
2 3 3
2 3 1
1 3
5 3 1 3 0 2
3 3 0 2
2 3 3
1 3
6 3 0 2 3 0 0
2 3 3
3 3 0 3
3 3 1 3
6 3 1 1 1 3 0
5 3 0 3 1 3
5 3 3 0 0 0
9 3 0 3 0 1 3 3 1 2
31 3 3 0 1 0 0 0 2 1 3 0 2 3 2 0 1 2 2 0 3 0 3 1 0 1 2 3 0 3 1 0
6 3 0 2 1 1 3
17 3 0 3 0 3 0 1 3 3 0 3 1 0 1 2 1 3
3 3 0 3
3 3 0 3
5 3 1 3 0 0
3 3 0 1
1 3
4 3 1 3 0
23 3 2 0 3 0 2 0 3 0 3 0 1 3 3 1 2 2 0 3 0 1 3 0
12 3 0 3 0 1 3 3 3 1 3 0 3
2 3 3
5 3 3 3 0 0
6 3 3 2 0 3 0
1 3
2 3 3
8 3 0 1 3 3 3 0 2
1 3
9 3 3 0 2 2 0 0 3 0
4 3 1 1 0
2 3 3
8 3 1 3 0 2 2 0 3
2 3 3
4 3 3 0 0
3 3 0 3
15 3 3 1 3 3 3 0 2 0 0 0 1 3 3 0
2 3 3
10 3 3 2 3 0 3 0 1 2 3
4 3 3 1 0
2 3 3
20 3 3 1 0 2 0 3 0 3 1 2 2 0 0 0 1 3 1 0 3
16 3 3 1 3 3 1 2 1 1 1 1 2 0 0 2 0
5 3 0 3 1 3
3 3 0 3
11 3 0 3 0 1 1 1 3 0 3 3
1 3
13 3 1 3 1 3 1 3 3 2 0 1 2 1
15 3 0 3 0 2 3 3 3 0 1 1 1 2 0 3
4 3 1 1 3
4 3 2 0 3
13 3 0 3 0 1 3 3 0 3 0 1 0 0
5 3 2 0 0 3
5 3 3 0 1 0
5 3 3 1 3 3
3 3 0 3
4 3 3 0 0
7 3 0 3 0 3 0 2
20 3 0 3 0 1 2 1 2 3 1 3 3 1 2 1 0 3 3 0 3
3 3 3 0
3 3 3 0
17 3 0 3 0 0 3 0 1 2 1 1 0 0 1 3 3 0
14 3 3 0 0 3 0 0 1 3 1 3 2 1 0
3 3 0 3
3 3 0 3
2 3 3
5 3 3 3 0 0
6 3 0 3 1 3 3
3 3 3 0
5 3 1 3 3 3
7 3 0 3 1 3 0 0
5 3 1 3 3 0
3 3 0 3
28 3 3 1 3 3 0 1 2 2 0 3 0 0 0 3 3 3 3 0 1 2 0 3 1 0 1 3 3
5 3 0 3 3 2
5 3 0 3 0 3
12 3 0 3 1 3 0 1 3 3 3 0 2
6 3 3 0 0 3 3
1 3
7 3 0 2 3 0 0 3
6 3 3 1 3 3 3
2 3 3
12 3 3 1 3 0 3 1 3 0 3 3 0
12 3 0 3 0 0 3 1 2 1 1 3 1
4 3 0 2 3
8 3 0 2 3 0 0 0 1
1 3
11 3 3 1 3 0 0 2 3 1 3 3
4 3 3 0 0
3 3 3 0
2 3 3
11 3 0 3 1 0 1 2 2 3 2 1
25 3 3 0 1 1 1 1 1 1 2 2 2 2 0 3 0 1 3 3 3 1 3 3 1 3
12 3 3 1 3 3 1 0 1 3 3 1 3
2 3 3
7 3 0 3 0 2 0 3
5 3 0 3 0 1
4 3 0 2 3
5 3 2 0 1 3
3 3 0 2
7 3 0 3 0 1 0 0
3 3 0 3
3 3 3 0
11 3 3 0 3 3 1 3 0 3 0 2
7 3 0 2 3 0 1 1
23 3 0 3 1 2 1 1 1 1 2 0 3 0 1 3 3 1 3 1 3 0 0 3
10 3 0 3 1 0 1 3 3 0 3
13 3 3 1 2 1 3 0 2 3 1 3 3 3
3 3 0 3
5 3 3 3 0 0
8 3 3 1 3 3 1 0 2
5 3 0 3 0 0
8 3 1 2 1 3 3 1 3
7 3 3 1 0 3 1 0
8 3 1 3 1 3 2 0 3
3 3 3 0
3 3 2 3
3 3 0 3
7 3 1 3 0 0 1 3
5 3 0 3 0 3
5 3 1 0 3 3
2 3 3
14 3 0 3 1 2 0 3 0 1 2 3 1 3 3
7 3 0 3 3 0 2 1
3 3 0 3
17 3 3 0 1 1 2 1 3 0 1 2 0 2 3 0 1 0
10 3 0 1 0 3 0 0 0 1 3
1 3
7 3 0 2 3 1 0 0
3 3 3 0
2 3 3
13 3 0 3 0 1 3 3 0 3 3 0 0 3
5 3 0 3 1 3
21 3 0 3 3 1 3 3 0 1 3 3 3 0 2 0 3 0 0 3 0 2
23 3 3 1 0 0 1 3 3 3 0 3 3 0 1 2 0 3 0 3 1 3 3 0
10 3 0 2 3 0 2 2 0 3 0
6 3 0 3 1 3 0
18 3 0 3 0 2 3 0 1 0 3 3 3 3 3 1 3 3 3
3 3 0 3
9 3 0 3 1 3 3 0 0 3
17 3 3 0 0 0 3 3 3 2 2 1 0 1 3 3 0 3
3 3 2 2
3 3 0 3
2 3 0
9 3 0 1 2 0 3 1 3 3
2 3 3
11 3 0 1 3 3 0 3 0 3 1 1
8 3 0 3 0 2 3 3 3
8 3 1 0 3 3 3 2 0
2 3 3
3 3 0 3
6 3 0 3 1 2 3
2 3 3
11 3 0 3 0 1 3 3 0 3 0 2
4 3 3 0 2
20 3 0 1 3 3 0 1 3 3 0 3 0 1 3 3 3 1 3 0 3
6 3 3 0 0 3 3
16 3 1 3 3 1 3 3 0 3 1 3 0 1 1 1 3
2 3 3
11 3 3 0 1 0 3 0 2 0 1 3
4 3 0 2 3
2 3 3
9 3 1 3 1 2 0 0 1 3
6 3 0 2 1 3 0
1 3
4 3 0 3 3
5 3 0 1 0 0
4 3 3 2 0
3 3 3 2
2 3 3
6 3 0 3 0 2 3
3 3 3 0
16 3 3 0 1 2 0 3 3 0 1 1 1 1 3 2 3
9 3 0 0 2 0 3 0 0 0
3 3 0 1
8 3 3 2 0 2 0 2 3
20 3 0 3 1 2 1 2 3 2 0 1 1 3 2 0 3 0 1 3 3
4 3 3 0 0
14 3 0 3 1 0 2 0 0 0 1 3 0 2 3
8 3 0 3 3 0 0 1 3
8 3 0 1 2 1 1 0 0
3 3 1 3
11 3 1 3 1 3 0 2 2 0 1 3
4 3 0 3 0
5 3 0 3 0 3
14 3 1 1 3 0 2 0 3 0 3 3 1 2 0
2 3 1
3 3 1 3
5 3 3 1 3 3
7 3 0 3 3 1 3 3
6 3 3 1 3 3 3
8 3 0 3 1 2 1 1 3
1 3
1 3
6 3 3 1 2 1 0
13 3 3 1 2 3 0 3 1 3 0 2 1 3
3 3 0 1
3 3 0 1
7 3 0 3 0 1 0 0
15 3 3 2 3 0 3 1 0 1 3 3 1 1 1 3
3 3 0 3
3 3 0 3
8 3 0 3 1 3 0 1 3
10 3 3 1 3 3 3 0 2 2 3
9 3 3 0 1 2 0 2 3 0
7 3 1 3 0 0 3 0
2 3 3
8 3 0 3 1 2 1 2 0
9 3 1 3 1 3 3 3 0 2
26 3 0 1 3 3 1 2 3 1 3 3 0 3 0 3 0 1 3 3 1 2 2 0 3 0 3
1 3
3 3 0 3
11 3 3 1 3 3 0 3 1 0 2 1
4 3 0 3 0
6 3 3 1 3 3 3
7 3 3 1 2 2 1 3
1 3
17 3 0 3 3 1 2 0 3 0 1 3 3 1 1 3 1 3
16 3 1 3 1 3 3 0 3 0 2 0 0 0 3 3 1
24 3 0 3 1 0 1 3 3 0 3 0 3 0 3 3 2 1 3 3 1 3 0 0 0
8 3 1 3 0 2 0 3 3
3 3 3 0
1 3
5 3 0 3 0 3
4 3 1 1 3
2 3 3
7 3 1 3 1 1 1 1
7 3 3 2 1 3 3 3
1 3
3 3 1 3
8 3 3 0 0 1 1 3 0
13 3 0 3 0 1 2 2 0 3 1 2 0 3
20 3 3 3 1 3 3 1 3 0 2 1 2 0 0 0 1 0 2 0 0
5 3 1 3 0 0
5 3 0 3 0 0
26 3 0 1 3 3 3 1 3 3 0 2 3 0 2 2 0 3 1 3 3 1 1 3 1 0 3
6 3 0 2 3 0 2
1 3
2 3 3
4 3 1 3 0
4 3 0 2 3
4 3 2 0 3
7 3 3 2 1 3 3 3
2 3 3
4 3 0 3 0
12 3 1 1 3 0 3 0 1 2 1 3 1
4 3 3 0 0
10 3 0 3 1 0 1 3 2 2 3
4 3 2 0 3
5 3 0 3 0 1
2 3 0
3 3 0 1
1 3
12 3 1 1 3 0 3 3 1 2 3 0 2
17 3 0 2 3 0 1 0 3 3 1 2 1 1 1 1 1 3
15 3 0 2 3 0 2 1 1 1 3 0 1 3 3 3
6 3 1 3 1 3 3
8 3 2 0 3 0 2 0 3
5 3 1 1 1 1
6 3 0 3 0 1 0
6 3 0 3 1 1 3
6 3 3 1 3 3 0
3 3 3 0
1 3
5 3 3 0 1 0
1 3
7 3 3 1 3 3 3 0
1 3
1 3
4 3 3 2 2
13 3 3 1 3 3 0 3 0 1 1 2 3 0
8 3 1 1 1 1 1 3 0
3 3 3 0
2 3 3
3 3 3 1
11 3 1 1 1 1 2 0 2 1 2 0
4 3 0 3 0
5 3 0 2 1 3
3 3 3 0
2 3 3
5 3 3 0 3 3
4 3 2 0 3
3 3 3 0
2 3 3
13 3 1 1 1 3 1 3 3 0 1 0 1 3
5 3 0 3 0 1
8 3 0 3 0 1 1 3 0
6 3 0 3 0 0 3
2 3 3
12 3 3 0 2 1 1 1 1 1 3 0 3
25 3 1 3 0 2 1 1 0 3 3 3 3 2 0 3 1 1 2 2 0 3 0 2 0 3
2 3 3
2 3 3
5 3 2 0 1 3
4 3 1 1 3
2 3 3
20 3 0 3 1 2 0 3 0 1 1 2 3 1 2 1 1 1 3 2 3
8 3 3 1 0 3 2 0 3
4 3 0 3 0
3 3 1 1
3 3 3 3
1 3
9 3 0 2 3 0 0 0 1 1
3 3 0 3
11 3 0 3 0 1 3 3 0 1 0 0
5 3 0 2 3 0
2 3 3
8 3 3 0 2 3 2 0 2
9 3 0 3 0 1 3 3 1 2
3 3 1 3
7 3 0 3 0 1 0 3
14 3 3 1 0 0 0 3 2 1 3 3 3 3 0
4 3 0 3 0
6 3 0 3 0 2 0
1 3
1 3
1 3
15 3 0 3 0 3 0 1 3 3 1 2 1 1 1 1
19 3 0 3 0 3 1 1 3 1 3 3 0 1 0 3 3 3 3 0
18 3 3 1 3 3 0 3 0 2 3 0 2 1 2 0 0 1 3
10 3 3 0 3 3 0 1 3 3 3
3 3 1 3
4 3 3 0 2
9 3 3 1 2 2 0 3 0 2
39 3 3 1 3 0 1 0 2 1 1 3 0 3 0 3 0 2 0 1 2 3 1 3 3 1 2 2 0 3 1 2 2 0 3 0 1 3 3 3
6 3 0 3 1 2 3
6 3 0 3 1 1 3
4 3 1 3 0
5 3 0 0 2 3
2 3 2
2 3 0
13 3 1 3 3 1 3 0 3 0 1 3 3 3
10 3 3 0 1 3 2 3 1 3 0
4 3 1 0 3
5 3 1 1 3 3
16 3 3 0 0 3 0 0 1 2 3 3 2 0 0 1 3
24 3 3 0 0 3 3 3 3 3 1 2 1 1 3 1 3 3 0 3 1 2 2 1 3
2 3 1
6 3 0 3 3 3 2
2 3 3
30 3 1 2 0 2 0 1 3 3 3 0 3 1 1 1 1 3 3 3 1 2 2 3 1 2 1 1 1 1 3
15 3 3 1 3 3 0 3 1 2 3 1 0 0 1 3
7 3 0 0 3 1 3 1
14 3 2 0 3 0 1 1 2 0 3 3 1 3 3
11 3 3 0 0 1 3 0 2 0 2 3
3 3 1 3
14 3 0 3 1 0 2 3 0 3 1 3 1 3 0
8 3 3 3 1 0 2 0 0
1 3
2 3 0
2 3 3
1 3
25 3 1 2 0 3 1 3 0 3 1 3 1 1 3 1 1 3 3 0 1 2 3 1 3 0
3 3 3 2
13 3 3 0 0 3 0 0 2 0 1 2 1 3
5 3 1 2 1 0
7 3 3 0 1 1 1 0
3 3 3 0
13 3 1 3 1 2 0 3 3 0 2 0 3 0
2 3 3
2 3 3
3 3 1 3
29 3 0 3 0 1 3 3 1 0 3 3 1 0 1 3 3 1 3 0 3 1 2 1 0 1 1 1 2 3
5 3 0 0 2 3
24 3 3 3 2 3 1 0 1 3 0 3 0 1 1 1 1 1 3 3 3 3 3 3 3
9 3 0 3 0 1 3 3 1 2
4 3 0 3 0
3 3 3 0
5 3 0 2 1 3
27 3 2 0 3 0 2 1 2 0 1 1 1 1 1 1 1 1 1 1 2 0 3 3 1 3 1 3
2 3 3
7 3 0 3 0 3 0 1
1 3
15 3 3 1 3 1 3 3 0 2 1 2 0 2 0 0
5 3 3 1 0 0
2 3 0
4 3 1 3 0
8 3 0 3 0 1 3 1 2
6 3 0 3 1 0 2
3 3 0 3
10 3 0 3 0 3 0 1 3 3 1
22 3 0 2 3 0 2 0 3 1 2 1 2 3 2 0 1 2 0 3 1 0 3
1 3
8 3 0 3 3 0 0 1 3
5 3 1 1 1 3
3 3 1 3
2 3 3
1 3
2 3 3
3 3 3 0
20 3 0 3 0 2 0 0 2 0 0 0 3 0 0 3 1 0 1 0 3
15 3 0 1 1 1 1 2 3 1 0 1 3 3 3 3
14 3 0 2 3 0 1 1 1 1 2 0 3 0 2
8 3 1 3 0 2 0 3 0
18 3 0 3 1 3 1 3 0 1 1 1 1 1 2 3 1 3 3
5 3 0 3 3 1
11 3 2 0 3 1 3 3 0 1 3 3
10 3 1 0 3 3 0 1 3 3 3
2 3 3
9 3 0 3 0 3 1 2 1 3
6 3 0 2 3 0 0
3 3 0 3
2 3 1
6 3 0 1 3 1 2
8 3 3 1 3 3 0 1 1
16 3 0 3 0 1 1 3 3 0 2 1 1 2 0 2 3
20 3 3 1 3 1 3 0 2 0 3 0 3 0 1 3 3 3 0 0 3
9 3 3 2 1 3 3 0 1 0
2 3 3
4 3 1 2 3
4 3 0 2 3
8 3 1 3 1 3 3 3 0
10 3 0 3 0 1 3 3 3 2 1
5 3 0 2 3 3
21 3 0 3 3 0 2 1 3 2 0 2 1 2 1 2 0 2 3 2 0 0
15 3 0 1 3 3 3 0 2 0 2 3 0 1 0 3
7 3 1 0 3 3 1 3
2 3 3
20 3 3 2 3 3 3 0 1 2 0 3 0 1 2 0 1 3 0 0 3
10 3 0 3 0 3 1 2 2 0 3
5 3 0 3 3 2
14 3 0 3 2 3 1 0 1 2 1 1 2 3 2
10 3 1 3 0 0 3 3 0 1 2
2 3 3
2 3 3
3 3 1 3
1 3
3 3 0 3
8 3 0 3 0 3 0 0 3
11 3 3 0 2 0 1 2 3 0 0 0
7 3 3 0 0 1 1 3
4 3 3 3 3
5 3 0 3 0 2
9 3 3 3 1 3 3 1 3 0
1 3
7 3 1 3 1 3 3 0
27 3 3 1 3 3 0 3 1 3 1 1 3 0 3 1 0 1 3 3 0 3 0 1 3 3 3 0
7 3 0 3 1 3 0 3
3 3 1 3
6 3 3 1 3 3 0
2 3 2
2 3 2
1 3
3 3 3 0
18 3 3 0 1 1 1 1 2 3 2 0 2 0 3 1 2 1 1
27 3 0 3 1 3 1 3 1 1 2 0 2 3 1 3 3 0 3 0 2 3 0 3 1 3 1 2
4 3 0 2 3
6 3 0 3 0 2 3
9 3 3 1 3 3 0 1 3 0
14 3 0 3 0 3 3 1 2 1 1 0 2 1 3
7 3 0 2 3 1 0 2
3 3 3 0
5 3 0 3 3 3
27 3 0 3 0 2 3 0 3 0 1 3 3 0 3 0 1 3 3 3 0 2 0 3 0 1 0 0
12 3 3 1 3 3 1 0 2 0 0 0 0
3 3 1 3
3 3 1 3
11 3 3 2 3 0 1 1 2 1 1 3
8 3 0 3 0 1 2 0 3
1 3
7 3 3 1 3 3 1 3
9 3 3 0 0 3 3 0 0 3
11 3 3 2 0 1 2 1 1 1 1 3
10 3 0 3 1 2 2 0 2 3 0
11 3 0 3 1 3 0 3 1 2 1 2
13 3 0 3 1 3 0 3 1 2 1 1 0 1
21 3 1 3 0 0 3 0 0 2 1 1 3 3 0 3 1 3 0 1 1 3
5 3 1 3 0 0
9 3 3 1 1 0 3 3 0 3
8 3 0 2 2 2 0 0 2
3 3 0 3
3 3 0 3
3 3 1 3
9 3 0 3 3 2 0 1 0 2
27 3 3 2 0 0 1 3 0 0 1 3 0 2 0 1 0 3 3 1 0 1 0 0 1 3 3 3
11 3 0 3 0 3 0 1 2 0 3 0
15 3 0 3 3 0 0 1 1 3 1 3 3 0 3 0
11 3 1 1 1 1 1 3 0 2 1 3
2 3 3
5 3 0 3 3 1
1 3
3 3 0 1
6 3 3 1 0 1 3
17 3 0 3 3 3 3 3 1 3 3 1 1 3 3 1 1 3
8 3 3 1 3 3 0 0 3
17 3 3 0 3 3 0 3 0 0 1 2 3 0 1 1 0 1
9 3 3 2 0 2 1 2 1 1
1 3
11 3 0 3 0 3 1 0 3 1 3 2
1 3
11 3 1 2 0 2 0 3 1 2 3 0
2 3 3
2 3 3
2 3 3
19 3 0 1 3 3 0 1 3 3 2 1 2 0 3 1 0 2 0 3
3 3 0 3
3 3 1 3
3 3 0 3
4 3 1 3 0
5 3 3 0 2 3
12 3 3 0 1 2 3 1 0 1 3 3 3
35 3 0 3 1 2 1 1 1 1 1 1 2 0 3 1 1 1 1 1 3 3 3 1 3 3 1 3 3 0 3 0 3 0 1 3
16 3 1 0 3 3 1 0 1 3 3 1 3 0 3 3 0
6 3 3 1 2 3 0
17 3 1 1 3 0 1 2 3 1 3 3 1 2 2 0 2 0
21 3 0 2 3 0 0 1 3 0 1 0 2 0 3 1 2 3 0 2 0 3
6 3 3 0 0 1 3
17 3 0 3 3 0 1 1 1 3 2 1 1 1 1 2 1 3
3 3 0 1
4 3 1 1 3
11 3 0 3 0 1 3 3 0 2 2 0
1 3
16 3 0 3 0 0 3 1 2 1 1 2 3 2 2 2 3
14 3 0 3 1 2 0 3 0 0 3 0 1 3 3
12 3 0 2 3 0 2 0 3 3 3 2 2
4 3 1 3 0
2 3 3
21 3 1 2 1 3 3 0 3 1 2 3 1 0 2 1 1 2 2 0 3 3
8 3 1 3 0 2 0 2 0
4 3 0 2 3
18 3 3 1 3 3 1 0 3 3 0 3 1 2 0 1 3 0 2
6 3 0 3 0 2 1
12 3 0 3 0 3 1 3 0 2 0 3 2
11 3 1 3 1 3 0 3 3 3 0 1
6 3 1 3 0 2 2
7 3 3 0 1 2 3 0
7 3 0 3 1 2 1 3
27 3 0 1 0 3 1 0 1 3 3 2 3 3 3 2 3 1 1 1 3 2 0 3 0 1 3 3
10 3 1 3 0 0 0 1 2 1 2
5 3 2 0 3 0
5 3 3 0 1 0
25 3 0 2 3 1 3 3 1 1 3 1 0 1 3 0 1 3 3 1 3 1 1 3 0 1
2 3 2
11 3 0 3 0 1 3 3 0 1 3 3
7 3 0 3 3 1 0 2
2 3 3
11 3 3 0 0 0 1 3 3 3 0 1
23 3 3 1 3 0 3 0 1 2 1 0 1 3 3 3 1 3 3 0 1 1 1 3
5 3 1 1 1 3
19 3 0 3 0 2 0 1 0 1 2 0 3 0 2 0 3 3 3 3
6 3 3 1 3 3 3
2 3 3
13 3 0 3 1 2 1 3 1 1 2 1 1 0
5 3 0 2 1 3
3 3 0 2
4 3 1 2 0
2 3 0
4 3 0 3 3
4 3 3 0 0
25 3 0 3 1 2 3 0 2 0 3 1 2 0 3 1 1 1 1 1 1 3 3 2 1 1
32 3 1 3 1 3 3 0 3 1 0 1 3 3 3 1 2 0 3 1 0 0 3 0 0 2 0 2 3 0 2 1 2
10 3 0 3 0 1 3 3 1 3 3
3 3 3 0
10 3 0 3 1 2 1 2 2 1 3
3 3 1 3
3 3 3 2
10 3 0 3 0 1 3 3 0 3 3
1 3
7 3 3 0 2 0 3 0
3 3 3 0
3 3 1 3
6 3 0 3 0 1 1
13 3 3 2 3 0 3 0 1 3 3 0 0 3
1 3
3 3 1 3
16 3 0 3 0 1 0 3 3 3 0 0 0 1 2 0 1
7 3 0 3 1 3 0 3
3 3 3 0
3 3 0 3
3 3 3 0
4 3 2 0 3
9 3 0 2 3 1 3 3 1 3
4 3 3 1 2
4 3 0 3 0
4 3 0 2 3
18 3 0 3 1 2 2 0 3 0 3 3 1 3 3 1 1 3 3
4 3 3 0 2
14 3 3 1 3 3 0 3 2 3 3 0 2 0 1
2 3 0
1 3
6 3 1 3 0 0 3
3 3 1 3
3 3 0 3
4 3 1 3 0
2 3 3
8 3 0 3 1 3 3 0 0
19 3 0 3 0 1 3 3 1 2 1 2 0 3 1 2 3 0 2 3
5 3 1 1 3 2
5 3 0 3 0 3
32 3 0 3 0 1 3 3 3 0 2 1 1 3 0 3 3 3 0 1 3 3 1 2 1 1 2 0 3 0 3 1 3
6 3 1 1 3 1 2
6 3 0 3 0 1 2
38 3 0 3 3 0 2 2 0 0 3 1 1 3 2 1 1 1 1 2 0 3 0 3 2 3 1 3 0 3 0 3 0 1 2 0 1 2 3
27 3 0 3 0 1 0 2 2 2 3 0 2 1 1 3 0 1 2 3 0 3 1 0 2 0 3 3
2 3 3
2 3 3
20 3 0 2 0 0 2 1 3 1 0 2 3 0 1 3 1 3 0 1 0
13 3 0 1 0 3 0 1 3 3 0 3 0 3
3 3 3 0
10 3 0 3 0 1 3 3 3 0 2
4 3 0 2 3
4 3 3 0 2
3 3 3 0
4 3 1 1 0
3 3 0 3
7 3 3 0 2 0 2 3
6 3 3 1 3 3 3
11 3 0 3 1 0 1 3 3 0 1 2
3 3 1 3
8 3 0 1 3 3 0 3 0
14 3 1 0 3 3 0 3 1 2 1 1 1 1 0
6 3 3 0 1 2 3
4 3 0 2 3
2 3 3
8 3 3 0 2 3 1 3 3
3 3 1 0
3 3 1 3
9 3 3 2 1 1 3 3 0 0
2 3 3
5 3 0 3 3 2
7 3 0 3 1 3 3 0
5 3 3 1 3 3
4 3 1 3 0
6 3 0 3 0 3 3
27 3 1 3 0 2 2 1 0 0 0 3 0 2 0 0 1 2 3 3 1 1 1 3 1 3 3 3
4 3 3 0 2
16 3 3 1 3 3 0 2 3 0 2 3 1 2 2 0 3
6 3 0 2 3 0 0
2 3 1
2 3 3
5 3 1 3 0 0
10 3 3 0 1 2 0 3 1 2 3
9 3 3 1 3 3 3 1 3 3
2 3 3
2 3 3
9 3 3 1 2 1 2 0 3 3
6 3 0 3 0 1 0
13 3 0 3 1 3 3 0 0 3 3 0 1 3
3 3 1 3
3 3 0 3
7 3 1 3 0 2 0 3
4 3 3 0 2
26 3 0 3 1 2 2 0 3 0 2 0 2 3 0 1 0 1 3 3 0 3 3 3 0 1 0
8 3 0 3 0 1 3 3 3
2 3 3
4 3 0 3 0
1 3
1 3
3 3 1 3
7 3 0 3 1 2 0 3
24 3 0 3 0 1 3 3 0 3 0 3 3 0 2 0 3 1 2 1 1 1 0 2 0
1 3
4 3 1 1 3
2 3 3
5 3 1 3 0 2
9 3 3 0 1 0 2 3 2 3
6 3 3 0 0 1 3
13 3 0 3 1 3 0 3 1 2 1 1 1 0
5 3 1 1 3 3
2 3 3
4 3 3 2 3
2 3 3
9 3 3 0 0 1 3 0 1 3
6 3 0 3 1 0 2
4 3 2 0 3
4 3 3 1 2
8 3 2 0 3 0 2 1 3
2 3 3
1 3
4 3 0 3 3
2 3 2
7 3 0 1 3 3 1 3
10 3 3 0 2 0 3 3 1 2 3
4 3 2 0 3
7 3 3 3 0 0 1 3
4 3 1 3 0
9 3 1 3 1 0 1 1 2 0
15 3 1 3 1 3 1 3 0 2 0 3 1 0 2 0
3 3 3 0
2 3 3
40 3 0 3 0 3 0 3 0 1 3 3 3 0 1 1 1 2 3 1 3 3 3 0 2 0 3 0 1 3 3 0 1 0 1 3 3 0 3 0 3
12 3 0 2 3 0 2 2 0 3 0 0 0
5 3 1 1 2 3
8 3 0 3 1 1 3 3 1
9 3 3 0 1 1 1 1 1 0
3 3 0 3
17 3 3 0 1 1 1 1 1 1 1 2 0 3 1 3 0 3
2 3 3
2 3 1
17 3 3 1 1 1 1 1 1 1 1 1 1 1 3 3 1 1
3 3 0 3
4 3 0 2 3
14 3 3 2 0 0 1 2 1 1 2 0 3 1 3
9 3 0 3 0 3 1 2 3 0
10 3 0 3 0 1 3 3 0 3 0
5 3 0 3 3 0
15 3 0 2 3 0 2 1 3 1 3 3 1 1 1 1
7 3 2 2 0 1 2 3
9 3 0 3 0 1 3 3 1 3
2 3 3
7 3 0 3 3 1 0 0
9 3 0 3 1 0 1 3 3 0
6 3 3 1 3 3 0
3 3 0 3
8 3 3 3 1 1 1 2 0
6 3 3 2 1 3 2
3 3 0 3
2 3 3
24 3 0 3 1 0 1 3 3 3 2 0 1 1 2 1 3 3 1 1 3 0 1 3 1
12 3 0 3 0 3 0 3 3 0 2 0 3
8 3 0 3 1 2 3 0 0
3 3 3 2
5 3 0 3 3 1
16 3 3 0 0 3 1 1 1 0 1 3 3 1 2 1 0
3 3 0 3
11 3 0 3 3 3 0 2 3 0 3 0
9 3 0 3 0 2 3 3 3 0
5 3 3 1 0 2
4 3 3 0 0
3 3 0 3
8 3 0 2 3 0 2 1 3
16 3 2 0 1 3 1 3 3 3 0 2 2 0 1 3 0
3 3 0 3
8 3 1 3 0 2 0 3 0
3 3 1 3
5 3 1 1 3 0
4 3 0 2 3
5 3 3 0 0 0
2 3 2
4 3 0 0 3
3 3 3 0
8 3 3 1 0 1 3 3 3
1 3
20 3 0 3 0 3 1 2 3 1 0 3 3 2 3 3 1 2 2 0 1
5 3 3 0 0 0
18 3 1 3 0 0 3 0 2 1 2 1 1 1 3 0 0 1 3
8 3 0 3 0 1 3 3 3
10 3 1 3 0 2 0 1 2 3 0
18 3 1 1 1 3 3 0 3 1 3 0 3 1 3 1 1 3 3
2 3 3
4 3 1 3 0
3 3 0 3
7 3 0 0 1 2 0 3
13 3 3 0 1 1 0 2 1 3 2 0 2 3
4 3 0 3 0
7 3 3 1 2 1 3 0
8 3 3 0 2 0 2 3 0
2 3 3
17 3 3 1 3 3 0 0 1 3 3 0 3 0 1 3 1 3
2 3 3
8 3 0 3 0 1 0 2 3
2 3 3
4 3 1 2 0
3 3 1 3
3 3 1 3
5 3 0 2 3 0
8 3 2 0 3 0 0 1 3
6 3 0 2 3 0 0
2 3 3
1 3
5 3 0 3 0 2
10 3 0 2 3 0 2 0 2 1 3
6 3 3 1 2 2 3
5 3 0 3 0 3
5 3 0 3 0 3
4 3 0 3 0
17 3 1 0 1 0 1 3 3 3 1 3 0 3 1 3 0 3
7 3 3 1 0 3 1 1
3 3 3 2
2 3 0
9 3 1 1 1 1 3 3 2 0
14 3 0 3 0 1 3 3 2 0 3 0 0 1 3
1 3
2 3 3
1 3
5 3 3 3 3 2
2 3 3
3 3 3 0
5 3 3 0 0 0
4 3 3 2 0
17 3 3 3 2 0 2 0 3 1 2 1 1 3 3 3 3 2
3 3 1 2
2 3 3
7 3 0 3 1 3 3 0
5 3 3 0 2 0
5 3 3 1 0 0
17 3 0 3 3 1 3 3 0 3 0 2 3 0 1 0 1 1
3 3 1 3
2 3 3
1 3
12 3 0 3 0 2 3 1 0 3 3 1 3
24 3 3 1 2 0 0 3 3 1 1 3 1 1 2 0 3 1 3 3 2 0 1 0 3
5 3 3 0 0 0
9 3 0 3 0 1 2 1 3 0
1 3
9 3 0 3 0 2 0 0 0 0
25 3 1 1 3 0 0 3 3 1 1 3 3 0 3 0 3 3 3 0 1 2 1 1 1 3
8 3 0 3 0 1 3 3 3
7 3 0 3 0 1 2 3
6 3 3 0 2 1 2
4 3 0 2 3
2 3 1
5 3 0 3 1 0
6 3 1 3 1 1 3
11 3 3 0 2 1 3 0 1 1 0 1
5 3 1 1 1 3
10 3 2 0 3 1 1 1 1 3 0
4 3 3 2 0
24 3 1 2 1 1 3 1 1 3 1 3 3 3 0 1 1 2 2 0 3 3 3 0 3
5 3 3 0 1 3
3 3 0 3
1 3
22 3 3 1 0 1 1 1 0 1 3 0 0 1 3 3 3 1 0 1 3 3 3
8 3 0 3 1 2 1 3 0
7 3 0 3 3 3 0 0
14 3 1 0 3 3 1 3 1 1 3 1 3 3 3
3 3 0 3
16 3 0 0 2 3 1 2 3 1 3 0 2 1 3 0 2
8 3 0 3 1 2 0 0 2
2 3 3
5 3 2 0 3 0
8 3 3 1 3 3 1 2 0
17 3 1 2 0 1 3 3 0 3 0 3 0 1 2 2 0 3
3 3 0 2
16 3 0 3 3 0 2 0 3 0 1 0 3 1 3 0 0
2 3 3
4 3 0 3 0
9 3 3 1 3 3 1 3 0 0
4 3 3 0 3
2 3 3
16 3 0 2 3 0 1 0 3 3 2 0 2 1 0 0 3
3 3 0 3
4 3 0 3 3
4 3 1 1 3
19 3 0 1 3 3 0 2 2 0 1 1 1 1 1 3 0 0 1 3
5 3 0 3 3 0
23 3 0 3 0 1 3 3 0 3 0 1 2 0 3 0 1 1 1 1 1 0 1 1
2 3 3
9 3 0 3 1 1 1 1 0 1
8 3 0 0 0 1 2 3 3
5 3 3 1 3 3
11 3 0 3 3 1 2 0 3 1 3 3
2 3 3
1 3
14 3 3 0 1 3 3 3 3 2 0 3 0 2 1
2 3 3
32 3 0 3 0 1 3 1 3 0 3 1 2 0 2 1 2 0 3 3 3 3 3 2 0 1 2 1 3 3 3 3 3
2 3 2
9 3 3 0 2 0 2 3 3 0
2 3 3
4 3 0 3 3
2 3 3
2 3 3
1 3
3 3 0 1
5 3 0 3 0 0
8 3 0 3 1 3 0 3 1
12 3 3 2 3 3 3 0 1 1 3 2 3
2 3 3
5 3 0 2 1 3
5 3 3 1 3 3
11 3 0 3 0 2 3 0 2 0 2 0
4 3 0 2 3
5 3 3 0 2 1
3 3 0 3
1 3
2 3 3
16 3 0 3 1 0 1 3 3 0 2 3 2 1 2 0 3
3 3 3 0
17 3 3 3 0 2 0 3 0 1 0 2 0 1 2 1 1 3
1 3
4 3 3 2 0
7 3 1 1 3 0 2 2
1 3
8 3 0 2 3 3 0 0 3
1 3
4 3 3 1 2
7 3 0 3 1 0 2 1
9 3 0 2 1 3 0 0 1 3
2 3 3
8 3 3 1 3 3 3 0 0
8 3 0 3 0 2 1 0 2
6 3 1 0 3 3 3
3 3 0 3
5 3 0 3 0 2
2 3 1
5 3 1 3 0 2
4 3 3 2 0
4 3 2 0 3
2 3 3
9 3 3 0 0 1 1 1 1 3
1 3
2 3 3
1 3
8 3 2 0 1 3 0 2 3
6 3 3 1 3 0 0
9 3 2 0 3 0 1 2 0 3
3 3 3 1
8 3 3 0 0 3 3 0 3
10 3 0 3 1 3 0 3 0 3 0
3 3 0 3
8 3 0 2 3 0 0 1 3
8 3 3 0 1 2 1 3 0
13 3 0 3 0 1 3 3 1 0 0 3 0 0
9 3 2 0 3 0 2 1 1 3
10 3 0 3 1 3 0 0 2 3 0
3 3 1 2
3 3 1 3
13 3 0 3 1 1 3 0 0 0 3 3 3 0
24 3 3 2 1 1 2 2 0 3 0 3 1 2 3 0 2 3 0 0 0 2 0 3 0
1 3
5 3 1 2 0 1
2 3 0
9 3 3 1 0 0 3 0 3 0
3 3 0 3
11 3 3 1 2 3 0 3 3 1 3 3
7 3 3 0 2 0 2 3
2 3 3
3 3 1 3
5 3 1 3 1 1
20 3 0 3 3 0 1 1 2 0 3 1 2 3 1 3 3 0 3 0 2
12 3 1 2 0 3 1 2 1 2 0 3 3
6 3 0 2 3 0 0
3 3 0 3
4 3 1 1 1
10 3 3 0 2 0 1 1 1 0 2
2 3 0
3 3 3 3
5 3 1 3 0 0
3 3 3 0
5 3 0 3 3 0
8 3 0 3 0 2 2 2 3
3 3 1 3
1 3
2 3 3
8 3 3 1 2 3 1 3 3
3 3 1 3
7 3 0 3 0 2 1 3
2 3 0
2 3 3
11 3 1 0 3 3 0 1 2 2 1 3
21 3 3 0 2 1 3 0 3 3 3 0 3 1 2 1 1 2 0 3 0 3
10 3 0 3 0 3 0 3 0 0 3
2 3 3
5 3 3 2 0 3
16 3 0 2 3 1 3 3 3 1 3 3 3 0 2 1 2
2 3 0
5 3 1 3 1 2
3 3 1 3
12 3 3 1 3 3 1 2 2 0 3 0 3
7 3 0 3 3 0 2 3
5 3 1 1 3 0
2 3 3
4 3 0 3 0
20 3 0 2 1 0 1 3 3 0 0 1 3 3 0 1 2 3 0 0 0
4 3 3 0 2
4 3 3 0 2
12 3 0 2 3 0 2 0 2 3 1 2 1
12 3 0 3 0 3 0 3 1 0 2 0 0
6 3 3 2 3 1 3
1 3
26 3 0 3 1 3 0 3 3 1 3 3 3 0 2 0 3 0 1 3 3 3 0 2 0 3 0
12 3 0 3 0 1 1 3 3 3 3 0 0
7 3 3 1 1 2 0 3
6 3 0 3 1 2 3
3 3 0 3
1 3
29 3 0 3 0 3 1 2 0 3 0 2 0 3 1 3 3 1 3 3 0 1 3 0 3 3 3 1 2 3
10 3 1 1 3 3 1 3 3 0 2
18 3 1 3 0 1 2 1 3 0 0 3 0 0 2 0 1 0 3
2 3 3
2 3 3
19 3 0 3 1 0 1 3 3 0 1 3 3 1 3 3 3 3 2 3
8 3 1 1 3 3 0 3 0
8 3 3 0 1 2 3 1 0
2 3 3
6 3 0 1 0 2 0
11 3 0 3 1 2 1 3 1 0 1 0
1 3
12 3 0 3 1 2 3 1 3 0 3 0 3
3 3 1 2
6 3 1 1 3 0 2
5 3 1 1 3 0
10 3 1 3 0 2 3 2 0 2 1
10 3 0 2 3 0 2 2 0 3 0
3 3 0 3
3 3 1 3
1 3
7 3 3 0 1 1 1 3
2 3 3
27 3 1 3 2 0 2 1 1 1 3 0 3 3 3 1 3 0 1 1 1 1 2 0 2 3 0 0
8 3 0 3 1 3 1 3 2
5 3 0 1 3 3
10 3 1 1 3 0 1 0 1 3 3
5 3 0 3 0 2
18 3 3 1 3 3 0 0 1 3 0 2 0 3 0 0 3 1 2
4 3 1 3 0
4 3 1 3 0
5 3 3 0 0 3
15 3 1 3 0 0 0 1 2 0 3 0 2 3 2 1
6 3 1 3 0 0 0
4 3 0 3 2
6 3 1 0 2 2 3
3 3 3 0
3 3 3 2
12 3 0 3 1 2 0 3 0 2 3 2 2
13 3 0 3 1 0 1 3 0 1 3 3 1 3
34 3 3 1 3 3 0 1 3 3 0 0 3 1 2 1 1 0 1 2 1 1 3 1 3 0 1 3 3 0 3 1 2 1 0
6 3 3 0 0 3 3
24 3 0 2 3 0 2 0 3 0 0 3 0 1 0 1 3 3 0 3 1 1 3 1 0
14 3 3 3 3 2 0 0 2 0 3 0 1 2 3
3 3 0 3
4 3 1 3 0
21 3 3 0 0 3 0 0 2 0 3 0 1 3 3 0 1 3 3 0 2 3
12 3 2 0 3 0 1 3 1 3 3 3 0
4 3 1 0 3
11 3 0 3 3 2 0 1 3 0 3 2
9 3 0 3 1 3 0 3 1 3
17 3 3 0 1 2 0 1 1 3 3 3 0 3 3 3 3 2
10 3 3 1 3 3 0 3 0 3 3
3 3 1 3
16 3 1 3 0 3 3 3 0 2 3 0 0 0 2 0 2
28 3 1 0 3 3 1 0 1 3 3 0 3 1 3 0 1 3 0 3 0 1 0 3 1 0 1 3 3
6 3 3 0 0 1 3
7 3 3 1 0 3 1 2
2 3 0
4 3 3 0 0
2 3 3
2 3 3
3 3 0 3
1 3
4 3 3 1 0
3 3 3 0
1 3
6 3 3 1 3 3 2
2 3 3
4 3 0 3 0
13 3 3 3 0 0 0 0 2 3 1 1 1 1
3 3 0 3
17 3 1 0 3 3 0 1 1 1 0 0 3 0 3 3 3 3
6 3 1 1 3 0 2
9 3 2 0 3 0 2 0 3 0
4 3 3 1 1
5 3 3 1 3 0
3 3 1 3
8 3 1 3 1 2 3 3 0
10 3 0 3 1 2 1 1 2 0 1
2 3 3
6 3 3 0 1 2 0
8 3 0 2 3 0 0 3 3
4 3 3 3 0
5 3 3 1 3 3
3 3 3 0
2 3 3
19 3 1 1 1 3 3 2 2 0 3 3 3 0 2 1 2 0 1 2
5 3 0 2 3 0
15 3 0 3 0 1 3 2 1 2 3 0 3 1 0 2
10 3 3 0 2 3 2 0 3 1 3
6 3 3 3 0 2 3
5 3 0 2 1 3
4 3 3 0 1
2 3 3
1 3
3 3 0 3
15 3 3 1 3 3 0 2 0 0 1 0 2 1 1 2
2 3 0
4 3 2 0 3
8 3 0 2 0 0 0 0 1
14 3 0 3 0 1 3 3 1 2 3 1 0 0 1
2 3 3
5 3 3 0 2 0
9 3 1 3 0 2 0 3 0 2
3 3 1 2
4 3 3 2 0
5 3 2 0 1 3
18 3 0 3 1 1 3 0 1 1 1 1 3 1 2 1 3 2 0
12 3 0 3 1 3 1 1 1 1 1 0 0
35 3 0 3 3 0 0 0 2 0 1 3 3 3 1 0 3 1 0 1 1 1 1 3 1 1 1 2 1 1 1 1 2 0 3 0
2 3 3
21 3 1 3 1 3 3 0 0 3 1 3 0 3 3 1 3 3 1 3 3 2
9 3 3 0 3 2 0 3 0 0
7 3 0 2 3 0 1 0
14 3 0 2 3 0 2 0 3 1 3 0 1 0 3
1 3
7 3 3 1 3 3 3 3
2 3 0
22 3 0 3 0 1 1 1 1 3 3 2 0 3 0 1 3 0 1 3 0 2 3
3 3 3 0
2 3 3
14 3 0 3 0 1 0 2 3 0 2 2 3 0 2
9 3 0 1 0 2 0 0 2 1
5 3 3 0 1 0
26 3 3 1 3 3 0 1 0 1 3 3 1 3 0 1 1 1 1 2 3 3 0 3 3 0 3
42 3 0 3 0 2 1 1 2 1 2 0 3 0 3 1 3 0 3 0 1 0 1 3 3 1 1 1 1 1 1 1 1 1 1 1 3 3 3 3 3 3 1
5 3 0 2 3 0
4 3 0 2 3
14 3 0 1 3 3 1 3 3 0 2 2 0 3 0
29 3 0 3 1 2 0 3 1 3 3 0 0 3 0 1 3 1 2 1 0 3 3 3 2 3 0 3 0 1
6 3 0 3 1 3 3
3 3 3 0
17 3 3 0 2 0 3 1 2 1 3 3 3 3 1 1 3 0
4 3 0 3 0
4 3 0 2 3
3 3 0 3
3 3 1 3
5 3 0 2 3 0
6 3 0 2 3 0 0
2 3 3
3 3 1 3
6 3 1 3 0 2 3
5 3 1 1 3 0
11 3 1 3 0 2 0 3 1 3 1 0
3 3 2 0
13 3 0 3 0 3 3 0 1 3 1 2 3 0
1 3
2 3 3
5 3 1 1 3 0
16 3 2 0 3 3 3 2 1 1 1 1 2 1 3 0 2
13 3 0 3 1 2 0 3 1 0 0 1 3 1
4 3 3 0 2
3 3 1 3
2 3 2
3 3 3 2
7 3 3 1 2 3 1 1
4 3 0 3 3
1 3
3 3 1 1
1 3
4 3 0 2 3
2 3 3
7 3 0 3 0 1 3 3
9 3 3 0 0 1 2 1 1 3
5 3 1 1 1 1
6 3 1 1 1 3 0
2 3 3
2 3 3
9 3 0 3 0 3 1 2 0 3
2 3 0
4 3 3 0 2
20 3 0 3 0 1 3 0 2 3 1 1 1 1 1 1 3 3 3 0 0
13 3 0 3 0 1 2 3 0 2 1 0 3 3
3 3 3 2
4 3 1 2 0
19 3 3 0 2 1 2 1 3 3 1 1 1 3 0 2 2 0 0 3
3 3 3 1
3 3 0 3
1 3
2 3 3
11 3 3 1 3 3 3 3 3 3 0 3
23 3 1 2 1 3 3 1 0 0 2 1 2 0 1 0 1 3 0 1 2 3 0 0
20 3 0 3 0 1 3 3 0 3 1 2 1 3 2 0 3 0 0 1 3
8 3 0 3 1 0 2 3 3
7 3 0 3 0 1 0 0
2 3 3
2 3 3
2 3 3
18 3 0 3 1 3 0 3 0 1 2 1 1 2 0 2 3 0 2
8 3 3 0 0 0 1 2 3
3 3 3 2
4 3 1 3 0
9 3 0 3 1 2 1 1 1 1
10 3 0 3 1 3 3 1 3 3 3
3 3 3 3
4 3 3 0 2
12 3 0 1 2 1 1 1 1 1 2 0 3
13 3 0 3 1 3 0 3 0 1 3 3 3 0
10 3 0 3 0 1 2 1 2 3 2
4 3 1 1 3
8 3 3 2 3 0 2 0 0
10 3 1 3 1 3 3 0 1 0 0
3 3 0 3
15 3 3 0 2 0 1 2 0 3 1 3 3 0 2 3
15 3 3 1 3 0 3 0 3 1 2 2 1 1 3 0
21 3 3 3 1 3 3 1 3 0 3 1 3 0 3 0 1 3 0 3 3 3
4 3 0 2 3
12 3 0 3 1 3 1 3 3 2 2 1 3
5 3 3 1 3 3
2 3 3
3 3 1 3
2 3 3
5 3 3 0 2 2
3 3 0 3
2 3 3
3 3 0 3
8 3 0 2 3 1 3 3 3
27 3 0 3 0 2 1 1 0 2 3 1 0 3 0 3 1 2 2 3 1 0 0 1 3 3 3 1
11 3 0 3 0 1 2 0 1 2 3 2
5 3 0 3 1 3
5 3 3 1 3 3
22 3 0 3 1 0 1 2 1 0 3 0 0 2 0 2 1 1 2 2 1 3 0
7 3 0 3 0 1 2 3
21 3 3 1 2 2 2 0 3 0 0 1 3 0 1 2 0 3 0 1 3 2
3 3 1 3
5 3 3 0 1 0
5 3 3 0 1 3
4 3 3 0 1
34 3 3 1 3 3 1 2 1 1 1 1 3 2 1 1 2 0 3 0 3 0 1 1 3 2 3 0 2 1 1 1 1 0 0
8 3 0 3 0 3 1 3 3
10 3 1 3 1 3 3 0 3 0 3
20 3 1 3 0 1 0 3 0 3 3 0 3 0 1 3 3 0 3 3 0
8 3 0 3 0 1 3 3 0
8 3 3 3 2 3 0 0 3
2 3 3
13 3 0 3 0 1 0 3 3 1 0 1 3 3
42 3 0 3 0 3 1 2 0 1 2 3 0 0 1 1 3 1 3 3 0 3 1 3 0 1 2 1 1 1 1 1 3 1 3 3 3 1 0 2 3 0 1
1 3
7 3 0 3 1 3 3 1
20 3 1 3 0 2 3 1 2 3 0 3 0 0 1 3 3 1 2 2 3
6 3 0 3 3 0 2
17 3 0 1 3 3 1 0 1 2 0 3 0 1 2 0 2 3
5 3 0 1 0 3
30 3 0 2 3 1 0 0 1 3 2 3 1 1 3 3 0 1 2 0 1 2 0 3 3 1 3 3 3 0 0
14 3 0 3 0 1 2 1 0 1 1 1 2 2 0
6 3 1 1 1 1 3
5 3 0 3 0 3
5 3 0 2 3 0
3 3 1 3
2 3 3
8 3 1 1 3 1 3 0 2
2 3 3
1 3
11 3 0 3 1 0 1 2 3 1 0 0
2 3 3
27 3 3 0 1 1 2 0 3 1 2 3 0 0 0 3 3 3 0 3 1 0 1 3 0 0 1 3
1 3
21 3 0 3 0 1 2 1 2 0 2 3 0 1 1 3 0 3 1 2 1 3
4 3 3 0 2
12 3 0 3 0 1 3 3 1 1 3 0 1
4 3 3 0 0
1 3
3 3 1 3
8 3 0 3 3 1 3 3 1
10 3 0 3 1 0 2 0 2 0 3
7 3 3 0 3 3 2 2
5 3 0 1 2 3
7 3 3 0 0 1 3 1
3 3 1 3
8 3 0 3 3 3 0 3 0
12 3 0 3 0 3 1 2 1 2 3 2 3
25 3 0 2 3 0 3 1 2 1 1 1 1 1 1 1 2 0 3 1 0 2 0 3 3 3
8 3 2 3 1 3 3 0 1
3 3 3 0
7 3 3 1 3 3 3 0
1 3
3 3 3 0
10 3 0 2 3 0 0 3 3 0 3
1 3
3 3 0 3
10 3 3 0 3 0 3 1 3 0 2
3 3 0 3
2 3 0
1 3
3 3 0 3
7 3 1 3 0 2 0 1
1 3
2 3 3
8 3 0 3 1 2 0 0 3
12 3 3 0 1 2 1 3 3 3 3 0 1
10 3 1 3 0 0 1 1 3 0 0
19 3 1 1 3 0 0 3 0 3 1 0 1 1 0 1 3 0 0 3
17 3 0 0 0 1 0 1 3 3 1 0 1 3 3 0 3 1
6 3 1 3 1 3 1
6 3 3 1 1 3 0
3 3 3 1
14 3 0 3 0 3 0 3 0 3 1 3 0 2 3
4 3 3 2 1
7 3 0 3 0 2 3 1
7 3 1 3 0 1 3 1
2 3 3
3 3 3 0
10 3 0 3 1 3 3 1 0 3 1
3 3 3 0
7 3 1 3 0 1 2 3
2 3 3
2 3 1
2 3 3
4 3 1 3 0
2 3 3
6 3 0 3 0 3 0
4 3 3 1 2
11 3 3 0 2 2 0 3 0 0 3 0
4 3 3 0 0
9 3 3 3 1 3 1 3 2 2
13 3 3 0 2 0 3 1 3 0 0 0 1 1
3 3 0 3
2 3 3
7 3 3 1 2 3 0 0
5 3 2 0 3 0
4 3 3 0 0
2 3 0
7 3 1 0 3 3 3 0
5 3 0 3 0 2
12 3 1 3 0 1 1 1 1 0 0 0 3
8 3 0 3 2 0 3 3 0
5 3 2 0 3 0
4 3 0 2 3
2 3 3
5 3 0 2 1 3
2 3 0
2 3 3
7 3 0 2 1 3 0 0
16 3 1 1 1 3 0 0 3 2 1 3 0 2 0 1 2
12 3 0 2 3 1 3 2 1 1 1 0 1
3 3 0 3
27 3 0 3 0 3 1 3 0 1 2 0 0 3 0 3 3 1 0 0 1 3 3 3 3 1 2 3
2 3 3
3 3 3 1
8 3 3 0 2 1 2 0 0
11 3 1 3 1 1 3 3 2 2 0 3
11 3 3 1 3 1 2 1 1 3 0 3
7 3 3 1 3 3 0 1
12 3 3 0 1 2 0 3 1 0 2 0 0
20 3 3 1 3 3 0 3 1 0 1 3 3 0 3 0 1 1 3 3 0
5 3 3 1 3 3
16 3 0 3 1 3 0 2 0 1 3 3 0 2 3 0 2
21 3 0 3 0 2 3 0 2 2 0 3 0 2 0 3 0 1 1 3 0 3
7 3 3 2 3 2 0 3
12 3 0 3 0 1 3 3 1 2 1 1 3
15 3 3 3 3 2 1 0 1 3 0 0 3 0 2 0
5 3 0 2 1 3
6 3 3 0 1 1 3
5 3 3 1 3 3
12 3 0 3 0 3 1 3 3 1 1 3 3
7 3 1 3 0 2 3 1
2 3 0
4 3 3 0 0
16 3 0 3 1 0 2 3 1 0 0 3 1 0 3 1 1
2 3 3
29 3 1 1 3 0 2 0 3 1 3 3 3 1 3 3 1 2 1 3 3 0 2 3 0 1 1 2 1 3
4 3 0 3 3
4 3 0 3 0
14 3 3 0 0 1 3 0 2 0 3 1 2 0 3
6 3 1 3 0 1 0
27 3 0 3 1 0 1 3 3 3 1 3 3 1 0 1 3 3 0 3 0 3 0 1 3 3 1 1
2 3 3
6 3 0 3 0 2 0
3 3 3 0
3 3 0 3
2 3 3
3 3 0 3
18 3 0 2 3 0 1 2 0 3 0 0 3 0 1 3 3 3 2
8 3 0 3 0 1 0 0 1
9 3 0 3 1 3 3 0 0 0
3 3 0 3
15 3 1 1 2 0 0 0 2 1 2 0 2 1 3 2
16 3 3 1 3 0 0 3 0 1 3 3 0 3 3 0 0
2 3 3
5 3 1 2 1 3
2 3 3
5 3 0 3 1 3
3 3 1 3
10 3 1 1 3 1 1 3 1 3 0
18 3 3 2 2 1 3 1 3 3 1 3 0 3 1 1 1 3 0
4 3 0 3 3
1 3
8 3 3 2 0 3 1 2 1
4 3 1 1 3
7 3 0 3 1 3 3 3
20 3 0 3 1 2 1 1 1 1 1 3 0 1 1 1 1 2 0 2 3
6 3 3 0 1 0 1
9 3 3 0 1 1 2 3 1 0
3 3 1 2
2 3 3
7 3 0 3 1 2 1 1
3 3 3 0
16 3 2 2 3 1 2 1 3 3 0 1 3 3 0 3 0
4 3 1 3 0
11 3 0 3 0 2 0 0 1 3 3 3
2 3 3
5 3 3 1 0 2
2 3 3
3 3 0 3
3 3 1 3
1 3
10 3 3 1 0 1 2 0 1 3 3
9 3 1 2 0 1 0 2 0 3
5 3 3 1 0 3
4 3 0 2 0
15 3 0 3 0 3 0 3 1 3 0 3 0 2 3 1
8 3 0 3 1 2 0 3 0
3 3 1 2
2 3 3
13 3 3 1 3 3 0 1 3 3 0 1 3 3
1 3
4 3 0 3 0
5 3 3 1 3 1
3 3 3 0
4 3 1 1 3
5 3 1 1 1 1
6 3 1 3 0 1 3
8 3 0 3 1 3 3 3 2
7 3 3 1 2 3 1 3
2 3 3
3 3 0 3
3 3 3 0
29 3 0 3 0 3 0 3 0 3 1 0 1 3 3 3 3 0 1 0 2 0 0 2 3 3 0 0 1 3
3 3 3 0
5 3 0 3 1 3
5 3 3 0 1 0
17 3 3 0 2 0 3 1 0 2 2 0 3 0 1 3 3 3
6 3 0 3 3 0 1
9 3 0 3 0 3 1 2 3 0
11 3 0 3 0 1 2 0 2 1 2 3
12 3 3 0 2 0 3 0 3 1 2 1 0
2 3 0
7 3 0 3 3 0 0 3
7 3 3 0 2 0 3 0
5 3 1 3 1 0
7 3 0 3 1 2 0 3
2 3 2
1 3
10 3 0 3 1 3 0 2 2 0 3
7 3 0 3 0 2 0 0
6 3 1 0 3 3 3
3 3 1 3
10 3 3 1 0 2 3 1 0 2 3
7 3 0 0 2 1 0 1
1 3
8 3 0 3 1 2 1 0 1
2 3 3
2 3 3
4 3 3 1 0
9 3 3 1 1 3 1 1 3 0
3 3 1 3
35 3 3 1 3 3 0 3 0 3 0 1 2 0 0 1 1 1 1 1 1 1 1 1 3 1 1 3 0 2 0 3 0 1 3 3
8 3 0 1 3 3 1 3 3
3 3 3 0
3 3 1 3
9 3 3 0 3 3 1 0 2 3
8 3 3 3 1 3 3 0 3
2 3 3
1 3
12 3 0 3 0 3 0 3 1 2 0 3 1
8 3 3 0 1 0 1 3 0
7 3 3 0 3 3 1 3
11 3 0 3 1 1 3 3 0 1 3 3
3 3 0 3
12 3 3 2 3 1 3 3 1 3 0 1 2
3 3 0 3
5 3 0 3 2 3
16 3 0 3 1 0 1 3 3 0 2 1 1 2 0 3 0
9 3 1 3 1 3 3 1 2 3
17 3 0 1 3 3 3 0 1 1 0 1 1 0 1 3 3 3
4 3 1 1 3
8 3 3 1 2 1 2 3 0
4 3 3 0 2
9 3 1 1 2 3 0 1 2 3
2 3 3
1 3
1 3
6 3 2 0 3 0 2
14 3 3 0 3 3 1 1 3 1 0 1 3 1 1
3 3 0 3
4 3 1 3 0
37 3 3 2 0 1 2 3 0 1 2 3 1 3 0 3 3 3 3 1 2 1 1 1 2 0 3 0 3 1 3 0 3 0 2 3 0 2
6 3 1 3 3 0 2
6 3 0 2 3 0 0
3 3 1 3
9 3 0 3 1 3 0 1 1 0
5 3 3 0 3 1
11 3 3 1 3 3 1 3 0 1 3 1
16 3 1 3 0 0 1 3 0 1 0 0 0 3 0 0 0
5 3 1 1 3 3
5 3 0 3 1 3
2 3 3
3 3 0 3
4 3 1 3 0
17 3 3 1 3 3 1 3 0 2 0 3 1 0 1 3 3 0
9 3 3 0 0 1 0 1 3 3
3 3 1 3
3 3 0 3
8 3 0 3 0 3 3 0 0
8 3 0 3 1 2 3 0 0
9 3 0 3 0 1 2 0 1 3
2 3 3
2 3 1
4 3 3 1 3
2 3 3
9 3 3 1 2 3 0 2 0 3
7 3 0 0 3 1 2 0
11 3 3 1 3 3 1 2 1 1 3 0
3 3 1 3
5 3 3 1 3 3
3 3 3 0
2 3 3
3 3 3 0
20 3 0 3 1 2 1 2 3 1 3 3 3 1 3 3 1 2 2 0 3
6 3 0 3 0 2 3
1 3
6 3 0 3 0 3 0
3 3 1 3
13 3 3 1 3 3 3 3 2 1 3 3 1 3
5 3 0 3 0 3
6 3 1 3 0 0 0
5 3 3 1 3 3
8 3 3 1 2 1 2 0 3
10 3 3 1 3 3 2 2 1 2 3
6 3 0 3 1 3 0
10 3 0 1 3 3 3 1 2 1 3
8 3 0 3 3 1 2 3 0
1 3
16 3 0 3 0 1 3 3 1 3 0 0 0 3 3 3 3
1 3
6 3 0 1 2 1 3
7 3 0 3 1 3 0 0
14 3 0 1 0 0 1 0 1 1 1 1 3 3 2
11 3 3 0 2 2 3 1 0 1 3 3
2 3 3
2 3 3
1 3
35 3 0 3 1 3 0 3 1 2 1 1 1 1 2 3 1 3 3 0 1 3 2 3 3 3 3 3 0 1 1 2 0 3 0 3
5 3 0 3 0 3
4 3 3 1 0
3 3 1 2
35 3 1 3 3 2 1 2 0 3 0 3 0 3 1 3 0 3 3 3 1 3 3 0 3 1 0 1 0 3 1 3 3 3 3 0
1 3
4 3 1 1 3
5 3 0 3 1 2
2 3 3
17 3 3 1 3 3 0 3 1 2 1 1 2 0 3 0 0 3
4 3 3 0 1
25 3 3 2 3 2 0 3 0 1 1 3 2 1 1 2 0 3 0 3 0 2 1 0 0 3
3 3 3 0
26 3 0 3 0 0 0 3 3 1 2 1 1 2 0 3 0 1 3 2 0 2 0 3 1 3 0
5 3 1 3 0 2
3 3 0 3
8 3 3 0 1 1 1 0 1
8 3 0 2 3 0 0 0 1
7 3 2 0 3 0 0 3
16 3 3 0 3 3 1 0 1 3 3 0 1 3 3 3 0
14 3 0 0 0 1 1 1 0 1 3 3 3 3 2
7 3 3 0 0 1 1 3
6 3 0 2 3 0 3
6 3 3 1 3 3 0
2 3 3
4 3 3 1 3
5 3 1 1 1 3
11 3 3 1 1 1 1 3 1 3 1 3
2 3 2
2 3 0
5 3 0 3 1 3
5 3 0 3 1 3
13 3 3 0 0 0 2 3 0 3 3 1 2 3
9 3 0 1 3 3 1 3 0 3
6 3 3 1 3 3 3
10 3 0 3 1 3 3 1 3 0 2
2 3 3
11 3 1 0 3 3 3 1 2 3 0 3
6 3 0 3 1 2 3
2 3 1
19 3 0 3 0 3 2 1 2 0 2 0 3 0 3 1 2 3 0 2
19 3 3 0 3 3 1 0 1 3 3 3 1 3 3 0 3 0 2 3
13 3 0 3 0 1 2 0 2 1 1 3 0 3
7 3 1 1 3 0 2 3
3 3 3 2
7 3 0 3 0 2 2 3
3 3 1 2
3 3 3 0
4 3 2 0 3
2 3 2
17 3 3 0 1 1 1 0 1 1 2 1 0 3 2 0 3 0
6 3 0 3 1 3 0
7 3 3 1 3 3 1 3
2 3 0
3 3 0 3
12 3 0 3 0 1 3 3 3 1 3 3 3
12 3 0 3 1 2 2 0 3 0 1 3 1
1 3
5 3 3 0 1 0
4 3 0 3 0
7 3 3 0 3 3 0 3
3 3 1 3
3 3 0 3
1 3
6 3 0 3 1 3 3
3 3 0 1
13 3 0 3 0 1 2 3 0 2 0 3 1 3
3 3 0 3
19 3 3 1 3 3 0 1 2 3 3 1 1 1 1 1 1 1 1 3
4 3 0 3 3
12 3 3 0 2 2 0 3 0 0 3 3 1
5 3 1 3 0 2
2 3 2
8 3 0 3 1 3 0 2 3
25 3 0 3 0 2 3 2 0 3 0 2 0 3 0 2 0 1 3 0 1 2 3 0 0 0
5 3 0 3 1 3
2 3 3
8 3 0 3 3 0 0 0 1
5 3 0 3 1 0
11 3 1 3 0 2 1 1 1 0 1 3
11 3 0 3 3 0 0 1 3 0 0 3
3 3 0 3
10 3 1 2 3 0 0 3 3 0 3
11 3 0 3 1 2 1 1 1 3 2 3
11 3 0 3 0 2 3 0 2 3 2 3
5 3 3 0 3 3
42 3 0 3 0 3 0 3 3 1 3 1 2 2 0 1 3 0 2 0 3 0 1 3 3 3 0 2 0 1 3 3 0 1 2 3 3 1 3 3 0 1 2
5 3 2 0 0 3
3 3 0 3
4 3 1 3 0
5 3 0 3 1 3
2 3 3
3 3 3 0
4 3 0 3 3
4 3 3 0 2
8 3 3 0 0 1 3 0 0
5 3 0 2 3 0
12 3 0 1 3 3 0 1 1 2 3 0 2
4 3 0 3 0
3 3 0 2
5 3 3 2 3 0
3 3 0 2
24 3 0 3 1 3 0 3 3 1 2 2 0 3 0 3 1 2 2 0 3 0 1 0 0
1 3
2 3 3
1 3
4 3 0 3 0
21 3 0 3 0 1 3 3 0 3 3 3 0 3 1 2 1 1 1 0 0 2
9 3 3 0 1 0 1 3 3 3
26 3 0 3 0 1 2 3 0 2 3 1 0 0 0 1 1 2 3 1 1 1 1 1 1 1 3
13 3 1 3 1 3 3 3 2 1 0 2 0 3
12 3 0 1 3 3 0 3 0 1 3 3 0
5 3 0 3 0 3
7 3 3 1 3 3 1 0
31 3 0 0 1 1 0 1 3 0 1 3 3 0 1 3 3 3 0 0 0 3 3 3 0 0 3 1 2 2 3 2
3 3 1 3
17 3 0 3 0 0 3 1 2 1 1 1 1 2 0 2 3 0
2 3 3
7 3 3 1 3 3 1 3
16 3 1 1 3 3 0 0 1 2 2 2 3 0 1 3 3
24 3 0 3 0 0 2 3 2 3 0 1 2 0 1 1 1 3 0 1 2 3 0 1 0
10 3 0 3 0 3 1 2 0 3 1
3 3 0 1
3 3 3 0
8 3 2 0 3 0 2 1 1
7 3 1 3 0 2 3 2
14 3 0 2 3 0 2 1 1 3 3 0 3 3 3
6 3 2 0 3 0 0
2 3 3
1 3
5 3 0 2 3 3
2 3 3
8 3 0 3 1 3 1 3 0
2 3 3
4 3 0 3 0
3 3 1 3
3 3 3 3
9 3 0 3 1 0 1 2 3 1
9 3 1 1 3 1 3 0 0 3
3 3 1 2
6 3 0 3 0 0 3
3 3 3 2
5 3 0 2 1 3
7 3 0 2 1 1 1 3
13 3 1 2 1 3 3 0 2 0 3 1 2 3
4 3 1 3 0
3 3 0 3
6 3 3 0 2 3 1
22 3 1 1 3 1 3 1 3 3 0 3 1 2 1 2 0 2 3 0 2 0 2
17 3 0 3 1 0 1 2 1 3 2 1 2 0 1 2 0 3
1 3
9 3 1 1 1 3 0 2 0 3
4 3 1 3 0
1 3
3 3 1 0
28 3 1 1 3 3 0 3 3 0 0 3 3 1 3 0 3 3 3 1 0 2 1 1 2 0 2 3 0
8 3 3 0 2 0 3 1 3
19 3 0 3 0 1 3 3 1 3 0 1 1 1 2 0 1 2 1 0
21 3 0 3 0 3 1 2 1 2 1 3 0 1 3 0 1 2 1 3 0 2
8 3 3 1 3 0 2 0 3
3 3 3 0
12 3 0 3 3 1 3 0 2 0 2 1 3
2 3 3
6 3 1 0 3 3 0
4 3 0 3 0
2 3 3
7 3 1 1 1 3 0 0
3 3 3 0
9 3 3 1 3 3 3 0 0 0
5 3 0 1 2 1
22 3 3 0 1 2 0 1 2 1 1 3 0 3 3 3 1 2 1 2 0 2 3
23 3 0 3 1 2 2 0 3 1 3 0 2 3 0 2 2 0 3 3 1 3 0 2
11 3 0 3 1 3 0 3 0 3 3 3
13 3 0 3 1 2 0 3 0 1 1 1 2 0
7 3 1 3 0 2 1 1
15 3 1 3 1 3 3 1 3 3 0 1 1 1 1 0
7 3 0 3 2 0 3 0
2 3 3
10 3 0 3 3 0 0 3 3 3 0
14 3 0 3 0 3 0 1 0 2 3 3 3 0 2
1 3
1 3
3 3 1 3
2 3 3
4 3 0 3 0
12 3 0 3 1 2 2 0 3 1 2 1 0
2 3 3
9 3 0 3 1 0 1 3 3 2
5 3 3 2 1 3
7 3 0 1 2 2 3 2
14 3 0 3 0 3 0 1 3 3 1 1 3 0 3
7 3 0 3 0 1 0 2
10 3 0 2 0 2 0 3 1 1 3
4 3 1 3 0
6 3 1 3 0 0 3
7 3 0 3 0 1 3 3
2 3 3
9 3 1 2 0 0 0 3 3 1
7 3 1 1 1 3 1 3
3 3 3 0
22 3 3 1 3 3 2 0 0 0 3 3 1 0 3 3 0 3 0 0 1 1 3
14 3 3 0 1 2 0 2 3 1 3 3 3 3 2
7 3 1 2 0 0 1 3
9 3 0 3 1 2 2 0 3 0
2 3 3
1 3
2 3 3
5 3 3 0 2 2
4 3 3 0 2
8 3 3 0 2 1 1 1 1
4 3 0 3 3
3 3 0 3
7 3 3 0 0 3 3 1
4 3 3 0 2
4 3 1 3 0
2 3 0
5 3 3 0 3 1
3 3 0 2
7 3 0 2 3 0 1 0
9 3 3 0 2 1 2 3 0 0
13 3 1 3 0 2 1 2 1 3 3 3 0 2
2 3 3
9 3 3 0 1 1 1 3 1 1
2 3 0
10 3 0 1 2 0 3 1 0 1 3
13 3 0 3 0 3 1 0 1 3 3 0 2 2
4 3 3 0 2
8 3 3 0 2 3 3 0 2
2 3 3
18 3 1 3 0 1 3 2 3 0 2 0 3 0 0 1 3 3 3
20 3 1 0 1 3 0 2 0 3 0 2 1 0 3 3 3 3 3 1 3
1 3
15 3 3 0 0 1 3 0 2 0 3 1 2 0 3 0
5 3 3 1 0 3
10 3 0 1 2 1 3 1 3 3 3
4 3 0 3 0
6 3 1 1 3 3 0
3 3 1 3
27 3 1 3 1 3 3 0 1 3 3 3 0 1 2 0 0 2 3 0 1 2 3 1 3 3 1 3
8 3 3 1 3 3 0 2 3
10 3 1 3 0 2 0 3 1 3 3
14 3 0 3 0 1 3 3 0 3 1 2 0 3 1
12 3 0 3 0 1 0 1 3 3 2 0 3
9 3 3 1 3 3 1 2 2 0
3 3 0 1
1 3
11 3 0 3 0 3 1 1 3 1 3 0
3 3 3 0
9 3 0 2 3 0 0 1 3 0
2 3 3
5 3 0 3 0 1
13 3 3 1 3 3 0 1 1 1 2 1 3 0
5 3 3 3 1 0
3 3 0 3
17 3 3 1 0 1 3 3 1 3 1 1 2 0 3 0 0 3
3 3 1 3
20 3 0 3 3 0 0 3 3 1 1 3 0 3 2 3 1 1 3 0 3
4 3 0 2 3
5 3 0 3 1 2
1 3
3 3 0 3
7 3 0 3 3 1 2 3
7 3 1 2 0 2 1 3
6 3 3 1 0 0 3
5 3 0 2 3 0
4 3 1 1 3
3 3 0 3
19 3 0 2 1 3 0 0 3 3 1 1 2 1 2 0 3 1 2 3
4 3 1 1 3
2 3 3
3 3 0 3
20 3 3 0 2 3 3 0 2 1 1 1 3 0 1 2 0 3 3 0 0
6 3 0 3 0 2 3
1 3
7 3 0 1 2 0 3 0
10 3 0 3 0 3 3 3 1 3 0
5 3 0 1 1 0
17 3 3 1 0 1 3 3 1 2 3 1 1 1 1 1 1 1
6 3 1 3 0 0 3
10 3 0 3 3 0 1 2 0 2 3
12 3 0 3 1 2 1 1 1 1 1 1 1
2 3 0
2 3 0
5 3 3 1 3 3
6 3 3 0 0 0 2
25 3 3 1 3 3 0 2 2 1 2 1 1 1 2 0 2 3 0 2 0 3 0 3 0 3
3 3 0 3
3 3 0 3
4 3 0 2 3
8 3 0 3 0 3 1 3 3
12 3 3 1 3 3 0 2 0 0 0 3 3
10 3 0 3 1 3 3 2 0 1 0
7 3 3 1 3 3 0 3
11 3 1 0 3 1 2 2 2 1 1 2
4 3 1 3 0
15 3 0 3 0 1 3 3 3 1 3 3 2 0 1 3
4 3 1 1 3
3 3 1 3
2 3 3
8 3 0 3 1 2 2 0 1
5 3 0 3 0 2
4 3 3 3 0
2 3 3
20 3 0 3 1 2 1 1 1 3 2 3 0 1 1 2 3 2 0 1 0
9 3 1 1 3 3 0 2 3 0
2 3 0
6 3 3 1 2 1 3
3 3 0 3
3 3 0 3
8 3 0 2 3 1 0 1 3
4 3 1 3 0
4 3 0 3 2
5 3 0 1 0 2
4 3 3 0 2
12 3 0 3 0 1 0 2 0 0 1 3 3
3 3 3 0
6 3 3 0 2 0 2
7 3 1 3 0 0 3 0
7 3 3 0 2 2 0 3
12 3 1 3 0 1 1 2 3 1 3 3 3
4 3 3 2 0
8 3 3 1 3 1 2 3 3
15 3 0 3 1 2 0 3 1 1 3 2 1 3 0 0
13 3 0 3 3 1 1 3 0 1 1 2 0 3
28 3 0 0 1 1 1 1 0 0 1 3 3 1 1 3 3 1 3 3 2 0 1 3 0 0 1 3 0
3 3 1 3
7 3 1 0 1 3 3 3
2 3 2
20 3 0 1 0 1 3 3 0 1 3 3 1 0 2 0 0 1 3 3 0
1 3
3 3 1 3
3 3 3 2
12 3 0 3 1 3 1 3 3 1 3 2 3
4 3 1 1 3
3 3 1 3
3 3 1 3
3 3 3 2
3 3 1 2
5 3 0 2 1 3
11 3 3 0 0 1 3 1 3 2 1 3
5 3 0 3 3 0
14 3 0 3 0 3 0 1 0 3 3 0 3 0 2
13 3 3 0 0 0 1 1 1 2 0 3 1 3
7 3 3 2 0 0 3 3
2 3 3
5 3 0 3 0 3
3 3 1 3
5 3 0 3 3 0
5 3 3 2 0 2
4 3 3 0 0
13 3 3 0 2 3 0 3 1 2 1 1 3 0
8 3 0 3 1 2 1 1 0
5 3 1 1 3 1
3 3 0 1
2 3 3
6 3 0 3 2 0 3
3 3 1 3
5 3 0 3 1 3
2 3 3
15 3 1 1 3 3 0 2 0 2 0 3 1 2 3 0
11 3 3 1 3 3 0 3 1 1 1 1
7 3 3 3 1 3 3 3
14 3 0 3 0 1 3 3 0 3 3 0 2 1 3
8 3 3 2 1 0 1 3 0
5 3 0 3 0 0
7 3 3 0 2 1 1 3
5 3 3 1 3 3
1 3
1 3
4 3 3 0 0
26 3 3 1 1 2 3 0 2 0 3 0 1 2 2 0 3 1 3 3 1 1 0 1 0 3 1
5 3 0 3 0 3
5 3 0 3 0 3
10 3 0 3 0 3 1 1 1 1 2
14 3 0 2 1 3 0 0 1 3 1 3 3 1 3
6 3 1 3 0 0 3
12 3 0 3 1 3 1 2 0 2 1 3 2
19 3 3 1 3 3 1 3 0 2 0 2 3 1 0 3 3 3 3 0
5 3 3 2 0 2
10 3 1 1 1 3 0 3 3 3 3
10 3 3 1 3 1 0 1 3 0 0
3 3 3 0
12 3 0 3 1 2 1 1 1 1 2 1 3
5 3 0 3 0 3
16 3 0 3 0 1 2 0 1 3 3 0 3 0 2 1 0
3 3 0 3
6 3 1 3 2 1 0
3 3 0 3
6 3 1 1 1 1 1
4 3 3 0 0
4 3 1 3 3
4 3 3 2 0
3 3 0 3
7 3 0 3 1 2 1 3
3 3 1 3
13 3 0 3 0 1 3 3 3 0 1 1 1 3
12 3 0 3 1 3 1 1 3 0 3 3 3
2 3 3
3 3 0 3
6 3 3 0 0 0 2
9 3 0 1 3 3 0 3 3 3
3 3 1 3
9 3 2 0 3 0 2 0 3 1
20 3 3 1 3 3 1 0 1 1 1 1 1 1 1 1 1 2 0 3 3
7 3 0 2 3 0 0 0
5 3 3 0 1 1
10 3 0 3 0 3 0 1 3 3 3
2 3 3
9 3 1 3 0 0 3 3 0 2
2 3 3
5 3 1 3 0 1
9 3 0 2 3 1 3 3 1 3
5 3 2 0 3 0
2 3 3
3 3 1 3
7 3 0 3 1 3 1 3
10 3 0 3 0 1 1 3 1 1 3
8 3 1 3 1 3 0 2 3
6 3 0 3 1 2 3
5 3 3 0 2 1
3 3 3 2
5 3 0 3 1 3
11 3 0 3 1 0 1 3 3 0 2 3
2 3 3
11 3 0 3 0 3 3 1 3 3 0 1
3 3 0 3
6 3 3 2 0 0 2
32 3 0 3 0 3 0 0 3 1 3 0 3 1 2 2 0 3 1 3 0 3 0 3 1 3 3 3 1 3 1 1 2
24 3 0 3 3 1 2 1 3 2 0 1 3 0 2 0 3 0 1 1 3 2 3 0 2
19 3 0 3 0 3 0 1 3 0 1 0 1 3 3 0 3 3 0 3
3 3 1 3
14 3 3 3 2 0 1 2 1 3 0 1 1 0 1
16 3 0 2 1 3 0 1 2 0 3 0 2 0 1 3 3
6 3 3 1 3 3 3
11 3 0 3 1 2 0 3 0 0 3 0
2 3 1
22 3 0 3 0 1 3 3 0 2 3 0 1 3 3 1 3 0 1 1 2 0 3
3 3 0 2
7 3 3 0 2 2 0 3
7 3 3 1 3 3 3 0
1 3
3 3 1 2
7 3 0 3 0 2 1 3
3 3 1 3
13 3 3 0 1 2 0 3 1 3 0 2 1 3
9 3 0 3 1 3 3 0 1 3
12 3 1 2 0 0 1 3 0 2 2 0 3
2 3 3
2 3 3
3 3 1 0
3 3 0 3
6 3 3 1 3 3 3
7 3 2 0 3 1 3 3
40 3 3 2 3 0 3 0 1 3 3 1 0 3 3 0 2 3 0 2 1 0 3 3 1 1 3 0 1 2 1 1 2 3 2 0 1 3 0 2 3
9 3 3 1 2 0 3 1 3 3
1 3
5 3 0 3 0 2
5 3 1 1 3 1
3 3 0 3
5 3 3 1 3 3
13 3 3 0 2 2 0 3 0 0 1 3 0 2
4 3 0 3 3
8 3 0 2 3 1 3 3 3
10 3 3 1 3 3 0 3 0 2 3
10 3 0 3 0 1 3 3 0 3 0
7 3 1 2 1 3 3 3
5 3 0 3 3 3
4 3 1 3 0
10 3 3 1 3 3 0 1 2 3 0
7 3 0 3 0 3 0 3
11 3 3 3 1 3 0 3 0 2 3 0
7 3 0 3 0 3 3 0
10 3 0 3 1 3 3 1 3 3 3
7 3 0 3 1 3 0 3
5 3 3 0 1 3
3 3 3 0
3 3 3 0
1 3
20 3 3 2 0 1 1 1 1 2 0 3 0 1 2 3 0 1 0 1 2
12 3 3 1 3 3 0 3 0 2 0 1 3
3 3 3 0
6 3 0 3 0 2 0
3 3 0 1
4 3 1 3 0
8 3 0 3 0 3 0 3 0
5 3 3 2 0 0
6 3 1 3 0 1 0
5 3 0 3 0 3
7 3 0 2 3 0 2 1
5 3 0 1 0 0
13 3 1 3 0 2 0 3 1 2 0 1 3 0
19 3 0 3 0 1 2 3 1 3 0 2 0 2 0 1 3 3 1 3
5 3 3 0 2 1
23 3 0 3 1 2 1 1 1 3 2 1 3 3 3 3 0 1 3 3 2 0 1 3
5 3 0 3 1 3
6 3 0 3 1 0 2
3 3 0 3
2 3 3
6 3 0 3 1 3 3
6 3 1 3 0 0 3
3 3 3 0
14 3 3 0 3 3 1 3 3 3 0 0 1 3 0
12 3 1 1 2 2 3 0 1 2 3 0 2
12 3 3 1 3 3 0 3 0 1 2 1 0
10 3 1 3 0 1 1 0 1 2 3
2 3 3
2 3 3
3 3 0 3
11 3 3 0 1 2 3 1 1 3 2 1
3 3 3 0
8 3 3 0 1 2 1 3 0
3 3 3 0
3 3 3 0
10 3 2 0 3 0 1 2 0 3 0
13 3 3 2 0 0 0 1 0 1 3 3 1 3
2 3 3
12 3 0 1 2 0 3 0 2 2 2 1 3
4 3 3 1 3
7 3 3 3 0 3 3 3
14 3 0 3 1 2 2 0 3 3 2 3 3 2 0
3 3 3 2
21 3 0 3 3 3 1 3 0 1 1 1 1 2 0 3 0 1 3 1 3 3
9 3 0 1 3 3 1 0 2 0
5 3 3 0 2 3
17 3 0 3 1 0 1 3 3 0 3 1 2 2 0 3 0 3
2 3 3
7 3 3 0 2 0 3 0
2 3 3
4 3 0 3 3
11 3 3 0 0 1 3 0 2 3 1 3
3 3 1 2
2 3 0
2 3 2
33 3 1 3 3 3 0 1 3 3 3 0 1 2 0 3 0 1 3 3 3 1 3 3 1 2 1 1 1 3 3 3 3 0
6 3 3 1 0 1 0
1 3
9 3 3 0 0 2 0 3 1 3
4 3 0 0 3
4 3 0 2 3
11 3 0 2 3 0 2 0 2 1 1 3
13 3 0 3 0 3 1 3 3 3 1 3 0 3
7 3 0 3 1 3 3 0
3 3 1 3
2 3 3
9 3 3 1 3 3 0 1 3 3
5 3 1 3 0 2
14 3 3 1 3 3 1 3 0 0 0 3 3 3 2
2 3 3
8 3 0 3 3 3 1 3 0
11 3 0 3 0 3 1 3 0 3 1 3
8 3 1 3 0 2 2 0 3
4 3 2 0 3
5 3 0 3 3 0
11 3 3 2 3 3 1 2 3 1 3 3
12 3 0 3 0 1 2 1 1 1 1 0 1
2 3 1
7 3 1 0 2 3 0 3
22 3 3 0 0 1 3 0 0 1 3 0 2 0 3 0 1 3 3 1 2 1 0
9 3 1 2 0 0 1 3 0 2
8 3 0 3 0 3 0 2 3
23 3 0 3 1 2 1 3 0 1 3 3 0 1 2 1 1 2 0 3 0 2 3 1
6 3 0 3 1 2 0
7 3 0 3 1 2 1 1
4 3 1 1 3
19 3 3 0 0 0 3 3 3 1 2 1 3 2 2 0 3 1 3 3
2 3 1
4 3 0 3 0
9 3 1 3 0 1 1 2 0 3
25 3 0 3 3 0 2 0 2 3 0 1 2 1 2 0 3 1 2 0 3 3 0 3 0 0
6 3 0 3 0 3 3
6 3 0 3 1 2 3
4 3 1 3 0
5 3 0 1 0 3
4 3 0 2 3
4 3 1 3 0
8 3 3 3 0 1 0 0 1
12 3 1 3 0 1 1 2 0 3 1 3 0
11 3 0 1 2 0 3 1 2 0 1 3
19 3 0 0 1 2 0 3 0 1 3 3 3 1 3 3 1 2 0 3
8 3 3 0 2 1 1 1 3
10 3 1 2 0 2 0 3 3 1 0
18 3 3 0 2 0 3 1 1 1 1 3 0 3 3 3 2 0 3
8 3 1 3 1 3 3 1 3
3 3 3 1
2 3 3
2 3 3
13 3 0 3 0 2 3 1 2 3 2 2 2 3
6 3 1 1 3 0 2
3 3 1 3
8 3 0 3 0 3 1 3 0
4 3 1 1 3
2 3 3
5 3 3 3 0 0
8 3 0 0 2 1 1 3 3
6 3 0 3 0 2 3
8 3 3 1 1 1 1 1 1
7 3 3 1 1 3 2 1
3 3 0 1
3 3 1 3
7 3 0 2 3 0 1 0
5 3 3 0 2 0
12 3 0 3 1 1 3 3 0 2 1 3 0
17 3 3 0 0 3 3 1 1 0 1 3 3 3 0 2 0 3
4 3 3 0 0
3 3 3 2
2 3 3
5 3 0 3 1 3
3 3 0 3
20 3 0 3 1 3 3 0 1 3 1 1 1 3 0 3 3 2 3 1 0
4 3 0 2 3
1 3
4 3 0 2 0
3 3 1 3
5 3 0 2 3 0
5 3 0 2 3 0
6 3 0 3 3 1 3
4 3 1 1 3
3 3 0 3
7 3 0 1 3 3 1 3
4 3 3 0 1
9 3 0 3 0 1 3 3 0 1
16 3 3 1 3 0 3 3 3 0 3 1 1 1 3 1 3
2 3 3
5 3 0 3 1 2
2 3 3
2 3 3
2 3 3
6 3 1 3 0 0 0
5 3 1 3 2 0
29 3 0 3 0 1 2 1 1 1 2 0 2 3 0 2 2 3 0 2 1 1 2 1 3 0 1 1 1 3
13 3 0 3 1 2 1 0 1 3 1 3 2 1
12 3 3 0 0 3 3 3 2 1 3 3 3
18 3 3 1 1 3 2 2 0 0 0 1 1 0 2 3 1 3 3
1 3
3 3 0 3
11 3 2 0 3 0 2 0 1 0 1 3
4 3 1 1 2
2 3 3
19 3 0 3 0 3 1 2 1 2 0 2 3 0 2 1 1 3 1 3
3 3 0 3
2 3 0
2 3 3
3 3 0 3
8 3 0 3 3 0 1 1 2
6 3 3 1 3 3 3
4 3 3 0 2
2 3 3
7 3 0 3 0 2 3 3
4 3 0 2 3
7 3 1 3 0 2 3 3
8 3 3 2 0 2 2 0 3
11 3 0 2 3 0 0 1 3 0 2 3
1 3
8 3 3 1 3 3 0 3 3
7 3 1 3 0 1 0 2
7 3 0 3 1 2 3 0
8 3 1 3 0 1 1 3 3
2 3 3
1 3
12 3 3 0 1 1 3 1 0 1 2 0 0
4 3 0 2 3
6 3 3 1 3 3 2
10 3 3 0 0 1 1 3 0 0 3
3 3 3 1
3 3 0 3
13 3 0 2 0 1 0 1 2 3 1 3 0 1
12 3 3 0 0 1 3 0 0 1 3 2 3
6 3 3 1 3 3 0
5 3 1 3 1 0
2 3 3
34 3 3 2 3 0 0 1 3 0 2 0 3 1 2 0 1 3 0 2 0 3 0 1 3 3 0 3 1 2 0 3 1 3 3
4 3 1 3 0
4 3 1 3 0
10 3 0 3 1 0 1 1 0 3 0
11 3 3 1 3 3 1 3 0 0 1 3
6 3 0 3 0 2 3
8 3 0 1 0 3 1 2 3
9 3 0 3 3 3 3 3 2 0
15 3 0 3 1 3 0 1 0 1 3 3 3 0 3 0
2 3 3
20 3 0 2 3 1 3 0 3 2 3 0 3 0 3 1 2 2 0 3 0
3 3 2 3
4 3 3 2 0
8 3 3 1 3 3 1 2 3
10 3 3 0 1 2 0 3 1 3 3
6 3 0 2 3 0 0
1 3
4 3 3 0 2
2 3 3
8 3 0 3 1 3 0 3 0
4 3 1 3 2
1 3
2 3 3
4 3 3 0 0
28 3 0 2 1 3 0 0 1 3 1 1 2 0 3 0 3 0 3 0 3 1 3 1 1 3 1 2 2
12 3 1 1 1 3 1 3 0 2 2 0 3
14 3 1 3 1 3 0 0 1 1 3 0 0 1 3
3 3 3 1
3 3 3 0
4 3 0 3 3
8 3 1 1 3 0 2 3 2
6 3 0 3 0 1 2
5 3 0 3 0 3
8 3 0 3 0 1 0 2 0
7 3 3 0 1 2 1 3
6 3 3 0 2 1 3
2 3 0
12 3 3 0 0 3 3 0 3 0 0 1 3
5 3 3 1 3 3
7 3 3 0 0 1 3 3
7 3 0 3 0 1 3 3
1 3
3 3 3 0
8 3 0 3 1 2 0 3 0
19 3 0 0 0 1 0 2 1 0 1 0 1 0 1 3 3 3 0 0
7 3 0 3 0 1 3 1
2 3 3
9 3 0 3 0 1 3 3 1 1
7 3 1 3 0 2 0 3
7 3 0 2 3 0 2 1
13 3 0 2 3 0 1 1 1 0 1 3 0 2
8 3 0 3 0 1 3 3 0
3 3 0 3
3 3 3 0
8 3 1 1 3 3 1 3 0
3 3 3 0
2 3 3
19 3 3 2 0 1 1 1 2 1 3 0 2 0 1 1 1 1 1 0
18 3 3 0 1 1 2 1 3 0 2 0 3 1 0 1 0 0 1
6 3 3 0 0 0 1
1 3
1 3
2 3 1
5 3 0 2 1 3
2 3 3
6 3 3 1 3 3 3
14 3 3 1 3 0 3 0 1 3 3 3 1 3 2
10 3 2 0 3 0 2 2 0 3 0
4 3 3 3 0
2 3 3
5 3 3 3 1 0
6 3 1 3 0 1 3
2 3 2
7 3 0 1 0 1 3 1
1 3
12 3 3 0 2 1 3 3 3 0 3 0 2
2 3 0
6 3 3 0 2 1 2
11 3 3 0 1 1 1 2 0 3 3 0
6 3 3 1 3 1 3
1 3
2 3 3
9 3 0 3 1 2 3 0 1 0
3 3 3 3
10 3 0 0 0 3 1 3 2 0 2
10 3 0 3 1 3 3 1 3 2 3
5 3 3 1 2 3
2 3 3
1 3
12 3 3 0 2 0 3 1 2 2 0 2 0
2 3 1
7 3 3 0 1 0 1 1
21 3 3 1 2 3 3 1 2 2 3 3 2 0 1 2 0 3 2 0 1 3
3 3 3 0
14 3 1 3 0 0 1 1 3 0 2 1 1 3 0
3 3 0 3
3 3 3 0
5 3 0 3 3 0
1 3
6 3 3 1 3 3 3
11 3 3 3 2 0 2 0 3 0 3 0
8 3 0 3 3 1 3 0 3
10 3 0 3 0 0 3 0 2 1 0
7 3 2 0 3 0 0 0
2 3 1
1 3
20 3 3 1 3 3 3 0 1 3 1 0 1 1 2 0 3 2 0 3 0
15 3 1 3 0 1 1 0 2 0 3 0 2 3 0 3
9 3 2 0 1 3 0 2 3 3
2 3 1
2 3 3
2 3 3
2 3 1
1 3
13 3 3 0 1 0 1 1 0 1 3 3 0 2
6 3 3 0 2 0 3
21 3 3 1 3 3 0 3 3 1 3 1 2 0 3 1 2 1 1 0 0 2
12 3 3 0 2 0 3 0 2 1 2 3 3
15 3 0 3 1 0 1 0 1 2 0 1 1 3 0 0
6 3 0 3 1 3 3
5 3 0 0 3 2
22 3 0 2 3 0 2 0 3 0 3 3 0 2 1 0 3 3 0 3 3 3 3
4 3 1 1 3
6 3 1 3 1 0 3
10 3 3 0 1 1 0 1 3 3 0
1 3
4 3 1 1 3
3 3 0 3
5 3 0 1 1 3
3 3 0 3
15 3 0 3 0 3 0 2 0 3 0 2 1 2 0 2
15 3 0 3 1 2 1 2 0 3 3 1 3 3 0 3
11 3 0 3 0 1 3 3 1 1 3 3
19 3 3 1 3 2 0 2 0 1 3 3 0 2 0 3 3 2 3 1
8 3 0 3 1 2 2 1 3
3 3 0 3
3 3 3 0
3 3 3 2
2 3 3
5 3 3 1 3 3
4 3 0 2 3
8 3 3 1 0 0 1 3 3
6 3 3 0 1 2 3
2 3 3
10 3 1 0 3 3 0 2 0 3 0
5 3 0 3 0 2
3 3 3 3
31 3 3 3 1 3 3 1 2 2 0 3 0 1 2 1 3 0 2 1 1 1 1 0 1 1 0 1 1 3 0 0
17 3 1 1 3 0 1 2 3 1 3 3 0 3 1 0 1 0
3 3 0 2
5 3 0 3 3 2
13 3 3 0 0 0 1 0 0 3 3 3 1 3
9 3 1 1 3 3 0 0 1 3
3 3 3 0
6 3 0 3 0 1 2
8 3 0 2 3 0 3 2 3
3 3 0 3
7 3 3 2 2 2 1 3
11 3 3 3 1 3 0 3 0 1 3 3
33 3 0 3 0 1 3 3 3 2 3 0 3 0 2 0 3 1 3 0 2 0 3 3 0 0 3 3 0 3 1 3 3 3
7 3 3 0 1 2 1 3
11 3 0 3 0 3 1 3 3 0 1 1
6 3 1 3 0 1 0
8 3 0 2 3 0 0 1 3
2 3 3
9 3 3 0 2 0 3 0 3 2
2 3 0
5 3 0 3 3 2
12 3 3 1 3 3 0 3 0 1 1 3 3
8 3 0 3 1 2 0 1 3
12 3 0 3 0 1 3 3 2 0 0 0 1
3 3 1 3
5 3 0 3 0 3
4 3 0 3 3
7 3 0 3 0 3 0 0
7 3 1 1 3 3 3 2
2 3 3
3 3 0 3
3 3 1 3
1 3
6 3 0 3 0 2 3
9 3 3 0 2 0 3 0 2 0
3 3 0 1
5 3 1 3 0 0
10 3 0 3 1 3 0 1 1 1 1
17 3 3 1 3 3 0 1 3 3 1 2 1 2 3 1 3 3
3 3 1 2
5 3 1 3 0 0
1 3
7 3 3 0 1 3 0 2
3 3 0 3
6 3 0 3 0 2 0
2 3 3
4 3 0 3 0
7 3 3 0 2 3 1 2
12 3 3 1 3 3 0 0 2 0 0 0 0
10 3 0 3 1 2 1 3 0 2 3
5 3 1 1 3 0
3 3 0 3
2 3 3
5 3 3 2 0 2
4 3 0 2 3
4 3 0 2 3
12 3 0 3 0 2 3 0 1 3 3 3 2
2 3 3
14 3 0 2 3 0 0 0 3 3 3 0 3 1 3
10 3 3 1 3 3 1 0 1 3 3
1 3
18 3 3 1 2 2 0 3 1 3 0 3 0 1 2 3 1 3 3
4 3 3 1 3
5 3 1 3 0 0
25 3 0 3 1 3 3 0 2 0 2 3 1 2 1 0 3 1 0 2 2 3 0 1 0 1
4 3 1 1 3
11 3 0 3 1 2 1 1 2 1 3 0
8 3 3 1 3 3 1 3 3
4 3 3 0 0
5 3 0 2 3 0
3 3 1 3
7 3 3 0 2 1 1 3
5 3 2 0 3 0
19 3 1 0 3 3 0 3 3 0 2 1 1 1 1 1 3 1 1 0
7 3 3 3 0 0 1 3
7 3 0 3 0 3 0 3
7 3 0 3 0 3 0 2
4 3 3 0 0
7 3 3 0 0 1 1 3
1 3
10 3 3 1 2 3 0 3 3 1 2
3 3 3 0
3 3 1 3
4 3 0 3 0
3 3 0 3
6 3 0 2 3 0 0
11 3 0 3 1 2 1 2 0 1 0 2
5 3 1 1 3 3
4 3 1 3 0
2 3 3
3 3 0 3
2 3 3
14 3 1 1 3 0 1 1 1 1 2 1 1 1 3
15 3 0 3 3 3 0 3 0 1 1 3 3 1 3 3
8 3 0 3 1 2 0 1 3
2 3 0
15 3 0 3 1 2 1 3 2 3 0 2 3 1 3 3
9 3 3 0 2 0 2 1 3 0
12 3 0 1 2 0 3 3 0 2 0 3 3
11 3 0 2 0 1 3 3 0 0 3 2
16 3 0 3 0 3 0 1 3 3 1 0 2 3 2 0 1
2 3 3
4 3 0 3 3
6 3 0 3 0 3 1
6 3 1 3 0 0 0
9 3 1 1 3 1 3 3 3 0
14 3 3 0 2 0 3 1 3 0 3 3 1 3 3
3 3 1 3
4 3 0 3 1
13 3 3 0 1 1 1 2 0 3 1 2 1 1
3 3 3 0
4 3 0 2 3
6 3 1 3 3 2 3
7 3 0 3 0 1 1 1
2 3 3
2 3 3
2 3 3
4 3 2 0 3
9 3 1 3 0 2 1 2 3 0
5 3 0 3 1 3
2 3 3
3 3 0 3
3 3 1 3
4 3 3 1 2
5 3 3 1 3 3
3 3 3 3
16 3 0 3 1 2 1 2 0 3 1 1 3 3 3 1 0
10 3 0 3 0 1 3 3 2 0 3
4 3 3 0 2
2 3 2
4 3 0 3 0
22 3 3 1 3 1 2 0 3 0 1 3 3 3 0 1 0 1 1 3 0 2 3
13 3 3 1 3 3 0 3 1 3 1 3 0 2
8 3 3 0 1 1 1 3 2
3 3 1 3
2 3 3
2 3 3
2 3 3
11 3 1 3 2 0 0 1 3 0 0 3
37 3 3 0 1 0 3 2 2 0 3 0 1 0 2 1 1 2 2 0 3 1 0 1 3 3 1 3 0 2 0 3 0 2 0 3 0 1
7 3 3 3 1 3 0 2
25 3 0 0 1 2 0 3 1 2 0 3 0 2 1 3 0 0 3 3 1 3 1 3 0 2
4 3 0 3 0
2 3 2
1 3
1 3
11 3 0 3 0 0 3 0 1 3 3 3
3 3 3 0
23 3 3 1 3 3 0 1 3 3 0 3 3 0 2 0 3 0 1 3 3 1 3 0
2 3 0
8 3 3 0 2 1 1 3 3
5 3 0 2 3 0
3 3 0 3
4 3 0 2 3
6 3 1 3 0 3 0
12 3 0 3 0 1 3 3 1 3 0 2 1
11 3 0 3 0 1 3 3 1 0 2 1
19 3 3 1 3 0 2 0 1 0 2 3 0 3 0 2 3 2 0 3
22 3 0 2 3 2 1 2 0 3 1 0 2 2 2 3 0 1 1 1 2 0 3
4 3 1 1 3
7 3 3 0 2 2 0 3
2 3 3
1 3
20 3 0 3 0 1 3 3 0 2 3 1 0 1 3 3 1 3 0 2 1
2 3 3
4 3 1 3 1
8 3 0 3 3 2 0 2 0
14 3 1 1 3 3 0 1 3 3 1 0 1 2 3
8 3 3 1 3 1 2 1 3
4 3 0 2 3
2 3 0
2 3 3
3 3 0 3
2 3 1
1 3
6 3 3 0 3 3 3
6 3 3 0 0 0 2
1 3
6 3 0 3 1 2 3
9 3 3 3 0 1 0 2 0 3
9 3 1 3 0 2 0 1 3 3
2 3 2
7 3 0 3 1 2 0 3
3 3 3 0
2 3 3
2 3 3
7 3 3 0 1 1 1 0
16 3 0 3 0 1 2 1 3 3 1 1 3 1 3 3 3
8 3 0 3 0 2 1 0 0
5 3 3 2 1 3
2 3 3
3 3 3 0
13 3 0 3 3 0 0 0 3 3 3 2 0 3
5 3 0 3 1 3
3 3 3 0
4 3 1 3 0
6 3 3 0 2 0 3
9 3 0 3 0 3 0 2 1 0
15 3 3 0 1 1 0 2 0 3 3 0 2 3 3 0
27 3 3 2 0 1 1 1 1 1 1 1 1 0 1 2 1 1 1 1 2 1 1 3 0 1 1 0
3 3 3 3
30 3 0 3 0 1 3 3 0 3 0 1 3 3 1 2 0 1 3 0 1 2 0 1 1 3 3 3 1 3 0
8 3 3 2 3 1 1 3 3
4 3 3 1 3
7 3 0 3 1 3 0 3
5 3 3 0 0 0
2 3 3
6 3 2 0 0 0 3
1 3
6 3 1 1 3 0 0
10 3 3 1 2 3 1 2 3 3 0
4 3 3 0 0
5 3 0 3 0 3
5 3 0 2 3 0
8 3 0 3 1 2 0 1 3
9 3 3 0 3 3 1 3 0 2
5 3 0 3 1 2
20 3 0 3 0 2 1 1 3 0 3 0 3 1 2 3 0 0 0 3 3
2 3 3
2 3 3
8 3 0 3 0 1 3 3 1
1 3
6 3 0 3 1 2 3
8 3 3 1 3 3 3 0 0
5 3 0 2 1 3
6 3 0 3 0 3 0
4 3 1 3 0
2 3 3
8 3 1 1 3 0 2 1 3
3 3 0 3
15 3 0 3 0 3 0 1 3 3 3 2 3 1 3 0
13 3 0 3 0 1 3 3 3 1 3 3 3 1
5 3 0 3 1 2
12 3 1 0 3 3 3 1 3 3 3 0 3
13 3 1 3 1 3 3 3 0 2 2 0 0 3
7 3 3 1 3 3 1 2
2 3 3
4 3 3 0 2
13 3 0 3 1 0 1 3 3 0 3 3 0 0
2 3 3
4 3 1 3 0
9 3 0 1 2 1 3 0 1 1
6 3 0 1 0 1 3
18 3 0 3 0 3 0 3 1 1 1 3 1 3 1 3 3 3 1
3 3 0 3
6 3 3 0 0 1 3
9 3 3 3 2 3 1 3 2 0
9 3 3 0 0 1 2 0 1 3
16 3 2 0 0 3 0 0 1 3 0 1 3 2 1 1 0
18 3 3 1 3 1 3 1 1 3 2 1 2 1 1 3 0 1 3
2 3 3
9 3 3 1 3 3 1 3 1 3
3 3 1 2
9 3 3 1 3 3 1 1 3 0
6 3 1 3 0 0 0
3 3 1 3
5 3 0 3 0 2
2 3 3
4 3 1 3 0
7 3 0 3 0 1 3 3
4 3 3 0 0
15 3 0 3 1 0 1 3 3 0 2 3 1 3 3 3
3 3 3 2
6 3 1 3 1 3 0
3 3 3 0
2 3 1
11 3 0 3 1 2 1 1 1 2 0 3
19 3 3 1 3 1 2 0 3 3 3 0 0 1 3 0 2 1 3 0
4 3 1 2 0
2 3 1
2 3 3
10 3 1 3 0 2 0 2 3 0 3
2 3 3
10 3 0 1 2 0 3 1 2 1 3
6 3 0 3 1 0 2
3 3 1 3
6 3 0 2 3 0 0
8 3 3 1 3 3 0 3 3
2 3 0
28 3 0 3 3 1 2 2 1 1 3 3 0 1 1 1 1 3 1 2 0 3 3 3 1 3 3 3 0
2 3 3
14 3 1 1 3 3 2 0 1 3 0 0 1 1 3
2 3 3
5 3 0 2 1 3
2 3 3
1 3
17 3 3 0 1 2 0 3 0 1 0 1 3 3 0 1 0 2
4 3 3 2 0
5 3 0 3 3 0
2 3 3
4 3 0 2 3
5 3 3 3 0 2
14 3 1 1 3 3 1 2 1 3 2 1 2 1 3
4 3 3 0 2
1 3
11 3 3 1 3 3 0 0 3 1 3 3
18 3 0 3 0 2 3 0 3 1 3 3 0 1 0 1 3 3 3
2 3 3
3 3 0 3
23 3 3 0 2 1 3 3 3 3 1 3 3 1 1 1 3 3 3 1 2 1 2 3
2 3 3
18 3 0 3 0 1 2 1 1 1 1 1 1 3 3 3 3 0 2
7 3 0 3 1 3 1 3
11 3 3 1 3 3 0 1 0 3 3 3
5 3 3 0 1 0
23 3 0 3 1 0 1 3 3 0 3 0 3 1 2 3 0 2 1 2 0 0 1 3
4 3 0 3 0
4 3 3 0 2
3 3 3 0
3 3 3 2
7 3 3 0 2 2 0 3
3 3 1 2
4 3 1 1 2
9 3 0 3 0 1 3 3 1 3
1 3
8 3 0 3 0 1 0 1 0
2 3 3
3 3 1 3
19 3 3 1 3 3 1 3 0 2 0 1 3 3 0 2 3 0 0 3
12 3 1 3 0 0 0 1 1 2 2 3 2
10 3 0 3 3 2 1 0 1 2 1
24 3 3 0 2 1 0 1 3 2 1 3 0 0 3 3 1 0 1 1 3 0 3 0 2
3 3 3 2
8 3 0 2 3 2 0 1 3
4 3 0 3 3
15 3 0 3 1 2 2 0 3 0 1 3 3 0 2 3
2 3 3
4 3 0 3 3
21 3 0 3 0 2 3 1 1 1 2 1 3 0 2 1 0 3 3 1 3 0
4 3 0 2 3
4 3 3 0 0
15 3 1 3 0 0 0 1 1 0 1 2 2 0 3 3
15 3 3 0 3 3 3 1 3 3 1 2 1 1 1 3
6 3 1 1 1 3 0
11 3 3 0 2 0 1 0 3 1 2 3
8 3 0 3 0 3 0 2 3
6 3 2 0 0 1 3
5 3 0 3 0 3
2 3 3
4 3 2 0 3
18 3 0 3 1 1 1 3 3 3 1 3 3 2 1 2 3 2 3
1 3
11 3 3 0 2 0 3 1 3 0 0 0
3 3 1 2
2 3 3
2 3 3
8 3 3 0 1 3 3 3 3
2 3 3
3 3 1 2
2 3 2
2 3 3
6 3 0 3 1 2 3
1 3
5 3 0 3 1 3
16 3 3 1 3 3 1 0 3 3 0 3 3 0 0 3 2
9 3 0 2 3 1 1 2 3 2
3 3 3 2
4 3 0 3 3
6 3 3 0 2 3 3
4 3 0 2 3
18 3 3 1 3 3 3 1 3 3 3 1 1 1 1 0 3 3 1
6 3 3 0 2 0 3
5 3 0 3 1 2
4 3 0 3 0
3 3 0 3
1 3
1 3
8 3 0 3 3 0 1 2 3
19 3 0 3 0 2 0 0 2 1 0 3 3 0 1 0 3 3 0 3
2 3 3
6 3 0 3 1 3 0
2 3 3
15 3 3 1 3 3 0 3 1 0 2 3 2 0 0 3
10 3 0 3 1 0 1 3 3 1 3
4 3 0 3 0
10 3 1 3 0 2 0 3 1 2 1
30 3 0 3 1 3 1 1 3 1 3 0 0 1 1 3 0 2 0 3 0 1 3 3 1 0 1 3 3 1 3
2 3 3
6 3 0 2 3 0 2
1 3
10 3 1 1 1 3 1 1 3 3 0
2 3 0
9 3 2 0 3 1 1 1 3 0
9 3 1 3 0 2 0 1 0 2
2 3 0
7 3 3 0 1 1 1 0
1 3
3 3 1 0
3 3 1 2
17 3 3 1 1 3 1 3 0 2 0 3 1 2 1 2 0 2
24 3 0 3 0 0 1 2 2 3 0 3 3 0 3 0 2 3 0 3 1 0 1 3 3
3 3 1 3
3 3 3 3
9 3 0 3 3 3 1 3 1 3
2 3 3
10 3 3 1 3 3 0 3 0 2 0
10 3 0 1 0 3 1 3 3 3 3
1 3
3 3 0 3
4 3 0 2 3
3 3 1 3
10 3 1 3 1 3 3 1 2 1 1
6 3 0 3 0 0 3
16 3 0 3 0 2 2 2 3 1 3 3 1 3 0 0 3
6 3 3 1 3 3 3
5 3 0 2 3 0
14 3 0 3 0 0 3 0 0 3 0 1 3 3 3
11 3 0 3 0 0 2 0 0 0 1 3
1 3
5 3 2 0 3 0
7 3 1 0 3 3 0 2
4 3 3 2 0
12 3 3 0 1 1 2 0 3 1 3 0 3
9 3 0 3 1 2 0 3 0 0
14 3 1 3 0 0 1 3 0 2 0 3 1 2 3
12 3 0 3 0 3 0 3 1 0 1 0 0
6 3 3 1 3 3 3
7 3 3 0 2 1 1 2
12 3 0 3 0 3 0 1 3 3 0 3 0
4 3 2 0 3
6 3 0 3 0 2 3
14 3 3 1 0 1 3 3 2 0 3 0 2 0 3
11 3 0 3 1 0 1 3 3 1 1 3
2 3 3
12 3 0 2 3 2 1 1 3 0 1 2 3
7 3 3 1 3 3 1 3
6 3 1 1 3 0 2
5 3 3 1 3 3
3 3 0 3
4 3 3 2 0
5 3 3 0 0 0
5 3 0 3 3 0
2 3 3
8 3 1 3 2 0 2 3 2
10 3 3 2 0 2 0 3 1 2 1
14 3 0 3 1 2 0 3 0 2 2 0 1 1 3
5 3 3 0 0 0
6 3 0 2 1 1 3
33 3 0 2 3 0 2 2 3 0 0 3 1 2 1 1 1 1 1 1 2 3 1 3 3 1 3 0 2 2 0 3 0 2
4 3 1 3 3
3 3 1 3
3 3 3 0
5 3 0 2 3 3
8 3 0 3 1 2 1 1 0
3 3 1 3
5 3 3 0 0 3
3 3 0 3
10 3 0 3 3 3 1 3 1 3 0
4 3 1 1 3
4 3 1 1 3
19 3 3 1 3 3 0 2 3 0 1 2 0 1 0 1 2 2 0 3
14 3 1 2 0 2 0 3 1 0 1 3 3 0 3
7 3 3 1 3 3 3 2
1 3
7 3 3 1 3 3 3 0
3 3 3 0
3 3 1 3
2 3 3
7 3 3 0 0 3 3 1
3 3 0 3
7 3 3 1 3 3 1 3
6 3 0 3 0 3 1
3 3 0 3
1 3
9 3 0 3 0 1 3 3 0 3
4 3 1 1 3
5 3 0 3 1 0
19 3 3 1 1 3 0 1 3 3 3 0 0 1 3 3 0 2 1 2
6 3 3 0 0 0 2
7 3 0 3 0 2 0 0
7 3 3 3 0 0 1 3
3 3 0 3
6 3 3 0 3 3 3
2 3 3
2 3 3
14 3 2 0 3 0 1 1 1 2 3 0 1 3 3
22 3 3 1 3 3 1 2 3 1 0 1 1 1 1 0 1 3 3 3 0 3 0
3 3 0 3
8 3 0 3 0 2 3 3 2
2 3 0
2 3 3
7 3 0 3 0 3 1 3
7 3 0 3 1 3 1 3
9 3 3 3 0 0 0 3 0 0
4 3 0 3 1
2 3 3
12 3 0 3 0 1 3 3 0 3 0 0 2
14 3 0 1 2 1 1 3 3 3 0 2 0 2 3
6 3 0 2 1 1 3
10 3 0 3 0 1 3 3 1 3 2
8 3 3 1 3 3 2 1 0
11 3 0 3 0 1 0 0 1 3 0 3
8 3 0 3 0 2 0 0 3
11 3 0 3 1 0 1 2 3 1 3 0
5 3 0 3 1 0
2 3 3
14 3 3 0 1 1 1 1 1 2 3 1 3 3 3
7 3 0 3 1 2 3 3
21 3 1 3 3 3 3 3 3 0 3 0 1 0 0 1 1 0 2 3 0 3
5 3 0 3 3 2
10 3 3 1 3 3 0 3 1 2 3
3 3 1 3
3 3 1 3
10 3 1 1 3 0 0 1 3 0 0
4 3 0 2 3
2 3 3
12 3 0 3 3 0 2 1 3 2 0 0 3
2 3 3
3 3 0 3
15 3 0 3 1 3 2 2 1 3 1 3 0 2 0 3
3 3 3 2
2 3 3
3 3 1 3
5 3 0 3 3 0
3 3 0 3
17 3 3 1 3 3 3 0 0 3 0 1 3 3 1 1 1 3
9 3 1 3 0 1 1 2 1 0
3 3 1 3
7 3 3 3 3 0 2 3
35 3 0 3 0 1 2 1 1 1 2 1 1 0 0 1 3 3 0 2 3 1 1 2 3 0 2 0 1 3 3 0 3 3 1 2
4 3 3 0 1
13 3 0 3 0 1 3 3 0 1 2 0 3 0
2 3 3
3 3 1 2
9 3 3 1 3 3 0 1 3 3
3 3 3 0
1 3
9 3 0 3 3 2 1 2 3 2
13 3 0 3 0 1 2 3 3 0 2 0 3 3
1 3
2 3 3
5 3 0 3 0 3
2 3 3
7 3 1 1 3 3 1 3
7 3 0 3 0 3 0 1
5 3 3 1 2 3
4 3 1 1 3
12 3 0 3 2 0 3 0 2 1 1 3 0
21 3 3 1 3 3 1 3 0 3 0 0 1 3 3 0 3 0 0 1 0 2
5 3 0 3 3 1
3 3 3 0
6 3 0 3 0 3 3
2 3 3
2 3 3
7 3 3 0 1 1 1 0
2 3 0
4 3 3 0 2
3 3 3 1
3 3 3 0
2 3 3
8 3 0 1 3 3 3 0 0
5 3 1 3 0 2
4 3 3 0 1
3 3 3 0
7 3 0 3 0 1 2 3
2 3 3
2 3 1
5 3 1 3 1 3
4 3 3 2 0
7 3 1 1 3 0 2 1
4 3 0 3 3
3 3 3 0
14 3 0 2 1 3 0 2 0 3 1 2 2 0 3
4 3 0 2 3
4 3 0 3 3
8 3 0 3 1 2 1 0 1
4 3 0 3 3
9 3 3 1 3 3 3 1 2 3
6 3 1 1 1 3 0
3 3 0 3
4 3 3 0 2
4 3 3 2 0
14 3 0 3 0 1 2 3 1 3 1 0 2 0 3
24 3 0 3 1 2 1 2 0 3 0 2 0 0 3 1 3 3 3 1 1 1 3 1 0
13 3 1 3 1 3 2 0 3 0 2 2 0 3
5 3 0 1 2 3
5 3 0 3 3 0
1 3
4 3 0 3 0
2 3 3
13 3 0 3 0 3 1 2 1 1 1 2 3 2
5 3 1 1 3 0
7 3 0 3 0 3 1 3
3 3 1 3
2 3 3
7 3 3 0 0 1 3 0
14 3 0 2 3 0 2 0 1 2 0 3 3 2 0
9 3 0 3 0 2 1 1 3 0
2 3 3
2 3 3
2 3 3
12 3 1 3 1 1 2 0 1 2 1 1 3
2 3 3
1 3
2 3 3
9 3 0 3 0 1 2 3 1 2
8 3 0 3 1 0 1 3 3
3 3 1 3
3 3 1 3
2 3 2
3 3 0 3
2 3 3
3 3 0 3
6 3 1 3 1 3 3
5 3 1 3 0 0
10 3 1 3 0 2 0 3 1 0 2
13 3 0 3 3 1 3 3 0 1 3 3 1 2
18 3 0 3 1 3 0 0 3 3 1 2 2 1 3 1 3 3 3
5 3 3 0 0 0
6 3 0 3 0 1 2
3 3 3 0
6 3 3 1 2 0 3
2 3 0
3 3 0 3
17 3 0 2 3 0 1 1 1 2 0 3 1 0 1 3 3 3
8 3 1 3 0 1 1 1 3
2 3 3
7 3 3 2 3 2 0 3
12 3 0 3 0 1 3 3 0 3 0 2 3
8 3 1 3 1 1 3 0 0
10 3 1 3 0 1 0 0 2 1 0
1 3
4 3 0 3 0
13 3 0 1 3 3 3 0 2 1 1 1 1 1
7 3 3 0 2 1 3 0
2 3 3
8 3 1 1 3 0 2 0 2
2 3 3
1 3
8 3 1 3 0 0 1 3 0
9 3 0 0 2 1 2 1 3 0
6 3 3 0 2 1 2
3 3 0 1
10 3 3 1 2 3 1 1 3 3 0
2 3 3
3 3 0 3
6 3 1 3 1 3 3
3 3 1 2
13 3 3 0 2 1 1 3 3 0 3 0 2 3
4 3 0 1 1
2 3 3
10 3 0 3 0 3 1 0 1 0 0
49 3 0 3 0 1 3 3 3 0 0 1 3 3 1 0 1 1 1 2 0 3 1 1 3 0 2 0 3 0 1 1 3 2 1 1 1 1 2 0 3 1 2 0 3 1 1 2 3 2
6 3 3 0 2 0 3
2 3 1
2 3 3
6 3 0 3 1 0 3
6 3 3 1 3 3 0
2 3 3
8 3 3 1 1 3 2 3 0
5 3 3 0 0 0
3 3 0 3
5 3 0 3 1 2
4 3 3 0 1
3 3 0 3
11 3 0 3 1 3 0 3 2 0 1 3
4 3 1 3 0
2 3 3
5 3 1 3 3 0
19 3 2 0 1 3 1 1 3 0 3 0 0 1 3 3 3 1 2 3
7 3 3 1 3 3 3 0
6 3 0 3 3 1 3
6 3 0 3 0 3 3
15 3 0 3 0 1 3 2 0 2 0 1 3 3 1 3
3 3 1 2
12 3 3 1 2 1 1 0 2 2 2 3 0
9 3 0 3 3 0 2 0 3 3
12 3 0 3 0 3 0 3 3 0 2 0 3
1 3
9 3 0 2 1 1 3 0 0 0
6 3 3 0 0 1 3
3 3 0 3
3 3 1 3
8 3 3 0 3 3 3 0 2
6 3 3 0 0 1 3
5 3 0 3 1 0
3 3 0 1
4 3 3 0 0
2 3 2
4 3 0 2 3
10 3 3 1 3 3 3 1 3 1 0
2 3 3
7 3 1 3 0 0 3 0
11 3 0 3 0 2 3 0 0 1 3 3
10 3 3 1 3 3 0 3 3 3 0
3 3 0 2
9 3 0 3 1 0 1 2 0 3
19 3 0 3 1 2 0 3 0 0 1 3 0 1 2 0 3 3 3 0
2 3 3
8 3 1 3 0 0 3 3 0
3 3 1 3
2 3 3
2 3 3
6 3 0 0 3 2 0
6 3 0 3 3 0 0
7 3 0 3 0 1 0 3
12 3 3 0 1 1 2 3 1 3 3 3 0
12 3 3 0 1 1 1 1 1 1 2 0 1
22 3 0 3 0 0 0 3 1 3 0 2 3 1 3 3 0 3 0 3 0 3 3
1 3
9 3 0 3 0 1 0 1 3 3
8 3 0 3 1 2 2 0 3
3 3 1 3
3 3 0 3
1 3
6 3 0 3 0 3 0
4 3 1 2 2
11 3 2 0 3 0 2 0 3 0 2 3
2 3 3
7 3 3 3 1 1 3 0
6 3 1 2 0 1 3
4 3 0 3 3
1 3
2 3 3
3 3 3 0
6 3 0 3 1 1 3
7 3 0 3 0 1 2 2
3 3 3 0
30 3 0 2 3 0 1 1 0 1 3 3 3 0 3 0 0 3 1 2 1 3 1 3 3 3 0 0 1 0 2
2 3 3
2 3 3
7 3 3 2 3 2 0 3
25 3 3 1 3 2 0 3 1 0 3 1 0 1 2 3 0 3 0 1 3 3 0 3 0 3
5 3 0 3 0 3
3 3 0 3
3 3 1 3
6 3 3 0 2 1 3
3 3 3 3
8 3 3 2 0 1 2 1 3
3 3 3 0
11 3 0 3 0 1 1 3 1 3 0 0
1 3
9 3 0 3 0 3 0 1 2 1
4 3 1 1 2
11 3 0 3 0 1 3 3 3 1 3 3
4 3 3 0 0
7 3 1 3 0 0 1 3
1 3
29 3 0 3 0 2 0 1 2 1 1 1 1 1 2 3 1 2 1 2 3 0 2 2 0 3 0 2 1 3
6 3 1 1 3 0 3
10 3 0 3 0 1 3 3 3 1 0
4 3 0 2 3
9 3 1 3 0 2 2 0 1 3
10 3 3 0 0 0 1 3 3 3 0
4 3 1 1 3
4 3 0 3 0
2 3 3
4 3 2 0 3
2 3 3
9 3 0 2 3 0 1 2 1 3
3 3 1 3
15 3 1 1 1 1 1 1 3 3 0 2 3 0 0 0
8 3 1 2 0 0 0 3 2
3 3 3 0
6 3 1 1 3 0 0
5 3 1 0 0 0
8 3 1 3 0 0 1 3 0
12 3 3 0 0 3 3 2 3 2 2 0 0
10 3 3 1 3 3 3 1 2 3 0
4 3 0 1 2
3 3 1 3
4 3 0 2 3
2 3 3
1 3
2 3 3
3 3 3 3
2 3 3
1 3
1 3
2 3 0
16 3 0 3 1 3 0 2 0 0 2 0 3 0 2 1 2
3 3 3 0
6 3 0 3 1 3 0
18 3 1 2 3 3 0 2 0 3 0 3 0 1 3 3 3 0 2
7 3 3 1 3 3 3 3
14 3 0 3 0 0 1 1 1 0 1 2 3 0 1
6 3 1 1 1 1 1
4 3 3 0 2
4 3 3 0 0
13 3 2 3 1 3 0 3 0 3 0 2 1 3
2 3 0
14 3 0 3 0 0 3 1 3 0 3 1 2 1 3
5 3 3 0 2 1
33 3 2 0 3 0 1 3 1 3 3 3 3 0 0 0 1 3 3 3 3 1 0 3 1 1 2 0 3 3 3 2 3 0
5 3 1 1 3 3
17 3 1 3 0 3 3 0 2 0 1 3 1 3 1 3 0 2
10 3 3 1 3 3 0 2 3 1 2
23 3 1 3 0 1 1 1 0 1 3 3 3 1 0 1 3 3 0 3 1 2 1 0
4 3 0 1 0
4 3 1 1 2
13 3 3 1 3 3 0 1 1 1 1 1 3 1
18 3 3 1 3 3 0 3 1 2 3 0 2 2 0 1 3 0 2
2 3 3
2 3 3
7 3 3 0 2 0 3 3
4 3 2 0 3
2 3 3
7 3 3 0 2 2 0 3
4 3 0 1 2
5 3 3 0 1 3
3 3 1 3
8 3 3 1 3 2 0 3 0
5 3 0 2 3 0
6 3 0 3 3 2 0
15 3 0 3 1 2 1 1 1 1 0 0 3 0 1 2
11 3 0 3 0 1 3 3 3 1 2 3
11 3 1 3 0 2 1 1 1 1 1 3
5 3 3 0 1 0
6 3 1 2 0 0 0
3 3 3 2
4 3 0 3 3
17 3 0 3 0 0 1 3 3 2 0 3 0 1 3 3 3 3
6 3 3 0 0 3 3
10 3 3 0 0 3 3 1 0 0 2
1 3
2 3 3
1 3
13 3 3 3 2 0 2 3 2 0 1 2 0 3
16 3 0 3 0 0 3 0 1 3 3 1 2 3 0 1 1
4 3 1 3 0
3 3 1 3
3 3 1 3
6 3 3 2 0 3 3
10 3 0 3 1 0 1 3 3 3 0
13 3 0 3 0 2 0 0 1 1 0 1 3 3
5 3 1 0 3 1
6 3 0 3 0 2 0
2 3 3
14 3 1 3 0 1 2 0 3 0 3 0 2 0 3
5 3 3 1 3 3
13 3 0 3 1 0 2 0 2 0 3 0 3 3
3 3 0 3
2 3 3
9 3 0 2 3 1 2 3 1 2
11 3 0 2 2 2 0 3 0 3 1 3
3 3 3 2
12 3 0 3 3 1 1 1 1 1 1 3 0
3 3 3 1
6 3 1 3 0 2 1
3 3 0 3
15 3 3 0 1 1 1 1 0 1 1 0 1 0 1 0
14 3 0 2 3 1 3 3 1 1 3 0 2 3 0
4 3 1 1 3
4 3 1 1 3
6 3 3 0 2 0 3
5 3 3 0 1 2
12 3 3 1 0 2 1 1 3 1 1 1 2
5 3 1 1 3 3
3 3 0 3
6 3 1 3 0 2 1
8 3 0 3 0 2 3 0 0
5 3 0 3 0 3
3 3 1 3
3 3 1 3
4 3 0 2 3
2 3 1
1 3
10 3 0 3 3 0 2 3 2 3 2
5 3 0 3 1 0
5 3 3 1 3 0
4 3 0 2 3
4 3 0 3 3
4 3 0 2 3
8 3 3 0 1 3 3 3 1
2 3 0
2 3 3
14 3 0 3 0 1 3 3 3 1 3 3 3 0 2
17 3 0 3 0 1 3 3 0 3 1 0 1 1 3 2 1 1
2 3 3
23 3 0 3 1 3 3 0 2 0 1 3 3 1 0 2 1 0 1 3 3 1 3 3
3 3 0 3
1 3
7 3 3 1 2 3 3 2
2 3 0
13 3 3 3 3 0 2 1 3 0 0 1 3 0
7 3 0 3 0 3 0 3
3 3 3 2
4 3 0 1 2
5 3 3 1 3 3
21 3 3 1 3 3 3 0 0 3 3 0 1 3 0 2 3 3 0 3 3 3
4 3 3 0 0
13 3 0 3 0 1 2 1 0 1 3 2 3 3
7 3 3 1 3 3 1 3
1 3
2 3 3
8 3 0 3 1 2 3 1 3
3 3 1 3
3 3 3 0
21 3 1 3 1 3 0 3 0 1 3 3 3 1 3 1 1 3 0 2 1 1
15 3 2 0 3 0 2 0 3 1 2 0 3 0 1 3
2 3 3
9 3 3 0 0 0 1 3 3 3
8 3 3 1 3 3 3 0 0
5 3 3 1 0 3
6 3 0 3 1 2 1
2 3 0
4 3 0 2 3
3 3 1 3
3 3 3 0
8 3 0 2 3 1 0 0 1
2 3 3
3 3 1 3
8 3 0 3 1 2 0 1 3
6 3 1 2 1 1 3
8 3 0 3 0 0 3 0 2
2 3 1
10 3 0 3 1 3 0 2 3 0 1
3 3 0 3
11 3 1 1 3 3 3 0 1 0 3 3
10 3 0 3 3 3 3 0 1 1 1
2 3 3
17 3 3 1 2 3 0 1 1 0 3 3 1 1 1 3 3 3
4 3 1 1 1
7 3 3 0 2 0 2 1
3 3 0 3
5 3 0 3 1 3
18 3 0 3 0 3 0 1 3 1 3 0 3 0 1 3 3 0 2
4 3 1 3 0
3 3 3 0
10 3 0 3 1 0 1 3 3 0 2
7 3 0 3 1 2 1 0
12 3 3 0 1 0 2 0 3 1 3 0 3
2 3 3
4 3 1 3 2
5 3 1 1 1 3
10 3 1 1 2 3 0 3 0 2 3
2 3 3
1 3
14 3 3 0 1 1 1 1 1 1 2 0 3 0 3
1 3
25 3 1 3 0 1 1 2 0 3 1 2 2 3 1 0 1 2 0 1 3 0 1 2 1 3
3 3 3 0
6 3 2 0 3 0 2
7 3 0 3 1 3 0 3
14 3 0 3 1 2 1 1 1 2 3 1 2 1 0
7 3 3 1 2 1 1 3
11 3 1 3 0 1 1 1 1 2 0 3
4 3 3 0 2
14 3 0 3 3 1 3 3 1 1 1 1 1 1 3
3 3 0 3
31 3 3 2 0 0 3 3 3 3 3 0 1 0 2 1 2 3 1 3 3 2 0 1 0 1 3 3 3 3 2 3
2 3 0
3 3 0 3
10 3 1 2 1 3 3 1 1 1 2
6 3 3 1 1 1 1
24 3 3 0 2 3 1 3 1 1 0 3 0 1 3 3 1 2 0 3 0 1 3 3 3
10 3 1 1 3 0 0 0 0 0 3
1 3
1 3
7 3 1 2 3 1 0 3
8 3 0 3 0 2 3 1 0
4 3 0 3 0
5 3 0 2 1 3
4 3 0 3 0
7 3 3 0 2 0 1 0
3 3 3 1
1 3
6 3 3 0 0 1 3
2 3 3
5 3 0 3 0 2
11 3 3 1 3 3 3 1 1 1 1 3
1 3
24 3 0 3 3 1 3 3 0 0 2 3 1 3 2 0 0 0 3 3 3 0 3 1 3
3 3 3 0
1 3
2 3 3
2 3 3
16 3 3 0 1 1 0 1 3 0 1 3 3 0 3 0 2
4 3 3 0 2
1 3
11 3 0 3 1 3 0 3 0 2 1 3
17 3 3 1 3 3 3 0 1 1 1 1 0 3 3 0 1 3
4 3 3 0 2
9 3 3 1 3 3 0 0 3 0
2 3 3
21 3 0 1 2 1 2 0 3 3 0 2 1 0 3 0 3 1 2 3 0 0
8 3 1 3 0 1 0 1 0
1 3
2 3 3
9 3 0 3 1 2 0 0 3 3
6 3 1 1 3 0 0
2 3 3
4 3 3 3 0
28 3 0 3 3 3 1 2 2 3 1 3 3 0 1 3 1 1 2 0 3 1 3 1 0 3 3 0 3
10 3 0 3 1 0 1 2 3 1 3
4 3 3 3 0
2 3 3
7 3 0 3 1 2 0 3
5 3 0 1 1 2
3 3 1 2
3 3 1 3
8 3 1 3 0 2 0 2 3
3 3 1 3
4 3 0 3 0
1 3
4 3 0 2 3
4 3 1 2 3
9 3 0 3 1 3 1 3 3 3
7 3 0 2 3 0 0 0
6 3 1 3 3 3 2
3 3 3 0
8 3 0 3 1 2 1 1 0
10 3 3 1 3 3 0 1 2 1 3
13 3 0 2 3 2 3 0 1 1 1 3 1 3
5 3 0 3 3 3
2 3 3
7 3 1 3 1 3 3 0
4 3 3 2 3
11 3 3 1 3 3 0 1 3 3 3 0
13 3 0 3 0 0 3 0 1 3 3 1 3 0
2 3 3
21 3 0 3 1 3 0 3 1 3 0 0 1 3 0 1 1 3 1 3 3 3
10 3 3 1 3 3 3 0 1 2 3
4 3 1 3 0
39 3 3 1 3 3 3 1 3 3 0 3 0 1 3 3 0 1 2 0 2 3 3 3 3 3 1 3 3 1 3 0 1 2 3 1 3 3 0 2
11 3 3 1 2 1 3 3 3 2 0 3
2 3 0
14 3 0 2 1 1 2 1 1 1 1 2 0 2 3
2 3 3
2 3 3
2 3 3
3 3 3 0
11 3 0 3 0 3 3 0 0 3 3 1
1 3
5 3 3 1 3 1
9 3 3 0 1 2 0 3 1 3
1 3
16 3 1 1 1 1 3 0 1 3 3 3 3 0 1 0 1
6 3 0 3 1 3 3
11 3 0 3 0 1 3 3 1 2 0 2
2 3 0
8 3 0 3 3 0 2 0 3
2 3 0
1 3
12 3 0 3 0 3 1 3 0 2 0 2 3
5 3 3 0 1 0
2 3 3
22 3 3 0 1 3 1 3 1 3 2 3 0 1 2 0 3 2 0 3 0 0 3
10 3 0 3 0 2 3 0 0 1 3
6 3 0 2 3 1 2
4 3 3 0 0
3 3 1 3
1 3
15 3 0 2 3 1 3 0 0 3 0 3 1 3 0 3
1 3
4 3 0 1 2
2 3 3
1 3
3 3 3 2
1 3
5 3 1 3 3 2
11 3 3 0 1 0 1 1 1 3 3 0
9 3 0 1 1 3 3 3 1 3
8 3 0 3 1 2 2 0 3
4 3 2 0 3
10 3 0 2 3 1 3 2 0 0 3
8 3 0 3 0 3 1 0 2
4 3 0 1 2
3 3 3 0
5 3 3 2 0 0
2 3 3
8 3 0 3 3 0 2 0 3
2 3 0
7 3 3 0 2 1 3 2
16 3 0 2 3 3 0 1 2 0 3 0 2 0 1 2 1
2 3 0
5 3 2 0 1 3
2 3 3
13 3 2 0 3 0 2 2 0 1 3 0 1 3
4 3 1 1 3
1 3
4 3 0 0 0
3 3 0 3
4 3 1 3 0
11 3 1 1 1 1 1 3 3 2 3 0
8 3 0 3 1 2 1 1 3
2 3 3
7 3 0 3 3 1 0 2
2 3 3
2 3 3
12 3 0 3 3 2 1 1 0 1 3 3 3
1 3
3 3 3 2
6 3 1 3 1 2 0
7 3 3 0 0 0 3 0
6 3 3 0 0 3 3
5 3 3 0 0 0
6 3 0 3 0 2 1
6 3 3 0 2 3 2
2 3 3
12 3 0 3 3 0 1 2 3 1 3 3 3
3 3 1 3
2 3 3
4 3 3 0 2
9 3 0 1 3 3 1 2 0 3
4 3 3 2 0
3 3 0 3
15 3 3 1 3 3 1 2 0 0 3 0 2 1 3 0
10 3 1 3 1 3 1 3 3 1 3
2 3 3
6 3 1 1 1 1 3
2 3 3
4 3 0 1 0
22 3 3 1 3 3 1 2 1 3 0 2 0 3 0 0 3 1 0 1 0 2 0
2 3 3
2 3 3
1 3
3 3 0 3
2 3 3
2 3 3
2 3 3
7 3 1 1 1 1 3 0
15 3 0 3 0 3 1 2 1 1 2 0 3 3 1 3
2 3 0
14 3 3 0 0 3 3 0 3 0 1 1 3 0 2
4 3 0 2 3
3 3 1 3
3 3 3 0
10 3 3 1 3 3 0 1 2 1 2
12 3 0 3 1 0 1 3 3 0 1 2 3
23 3 3 1 3 3 0 1 3 3 0 3 0 0 3 0 2 2 2 1 3 1 1 1
12 3 0 3 1 3 0 3 3 3 2 0 3
20 3 0 3 0 0 3 1 2 2 0 0 1 3 3 1 2 0 3 0 2
2 3 3
9 3 0 3 0 1 2 1 1 3
3 3 3 3
1 3
4 3 0 2 3
8 3 3 0 2 0 1 0 2
2 3 3
10 3 1 1 1 3 2 0 0 3 0
3 3 3 0
8 3 0 0 0 1 2 3 0
4 3 1 1 3
4 3 3 1 3
4 3 1 1 3
5 3 1 3 0 2
3 3 1 3
5 3 3 1 3 3
2 3 0
5 3 1 1 1 2
4 3 2 0 3
8 3 3 1 3 1 2 0 3
9 3 1 3 0 0 3 3 0 3
8 3 2 0 3 0 2 0 2
3 3 3 0
2 3 3
3 3 3 1
5 3 3 0 1 3
4 3 0 3 0
7 3 3 0 1 2 1 3
6 3 0 3 1 1 3
4 3 0 3 3
1 3
13 3 3 0 0 1 1 3 0 0 3 3 1 1
5 3 0 3 0 1
4 3 0 3 1
17 3 0 3 0 1 3 3 1 3 0 3 1 2 1 2 1 3
27 3 3 1 3 3 3 0 3 3 1 3 0 3 1 2 1 1 1 1 1 1 2 0 3 1 3 0
10 3 0 3 1 2 1 1 3 0 1
9 3 1 3 2 0 2 0 3 0
12 3 0 3 0 1 3 3 0 0 1 0 3
2 3 3
3 3 1 3
4 3 0 3 3
10 3 0 3 1 3 3 0 2 0 3
2 3 0
18 3 0 3 3 3 0 2 1 3 0 1 2 3 1 3 3 3 0
2 3 0
7 3 1 3 0 2 0 1
4 3 3 0 1
3 3 1 3
1 3
4 3 0 1 0
14 3 3 1 3 1 2 1 0 1 3 0 0 0 1
7 3 1 1 1 3 0 2
2 3 3
4 3 3 1 3
14 3 0 3 3 0 1 2 0 3 0 3 0 1 2
18 3 1 1 0 3 3 0 3 1 3 0 3 1 3 0 2 0 3
6 3 1 3 0 2 3
20 3 1 1 3 0 3 1 2 0 3 0 2 1 1 1 3 3 0 0 2
4 3 3 1 2
3 3 3 2
5 3 3 0 2 0
16 3 3 0 2 0 3 1 3 3 1 3 3 3 0 1 0
1 3
6 3 0 3 1 2 3
3 3 0 3
10 3 0 1 3 3 3 1 0 0 1
4 3 0 3 3
3 3 3 0
5 3 0 3 1 2
1 3
3 3 1 3
1 3
4 3 1 3 2
4 3 0 3 3
3 3 0 3
3 3 3 0
12 3 0 2 0 1 2 0 3 0 0 0 1
17 3 0 1 2 1 2 0 3 3 0 2 0 3 1 2 0 3
2 3 3
2 3 3
2 3 3
4 3 3 3 3
7 3 3 1 3 3 0 1
3 3 0 3
14 3 1 3 0 2 0 3 0 1 3 3 1 3 0
12 3 3 0 0 1 3 1 1 1 1 1 3
4 3 0 3 0
33 3 3 0 1 1 3 3 3 1 1 3 1 3 0 0 0 2 1 3 0 1 1 1 1 1 0 1 3 3 3 1 2 2
3 3 0 3
14 3 3 1 3 1 3 1 1 1 1 3 3 0 2
33 3 0 2 1 1 3 0 2 1 1 3 1 3 0 0 3 3 3 3 3 1 1 1 1 3 3 0 0 1 2 3 0 2
12 3 0 3 1 2 0 1 1 3 0 0 0
2 3 0
10 3 3 1 1 1 0 3 2 2 3
7 3 0 3 0 1 0 0
5 3 3 0 1 0
3 3 0 3
14 3 0 1 3 3 0 1 2 3 3 0 2 0 3
2 3 3
2 3 3
7 3 0 3 2 0 3 3
4 3 0 2 3
6 3 1 3 0 0 3
5 3 3 0 1 3
12 3 0 1 1 2 3 1 0 0 3 0 3
3 3 0 3
9 3 0 3 0 1 3 3 1 3
4 3 0 3 0
5 3 0 3 0 3
6 3 0 3 3 0 1
13 3 3 1 3 3 0 2 3 2 0 1 1 3
2 3 3
22 3 0 3 1 2 1 2 0 3 1 0 2 1 3 0 1 1 1 3 2 0 3
2 3 2
3 3 1 1
26 3 0 1 3 3 1 3 0 0 1 3 1 3 3 1 3 0 3 1 2 3 0 1 2 0 3
9 3 0 3 0 1 2 3 0 3
2 3 2
2 3 0
1 3
21 3 0 3 0 1 3 3 0 3 1 2 1 1 2 0 3 1 2 0 3 0
10 3 0 3 0 1 1 3 3 1 3
15 3 0 1 2 2 0 3 0 1 1 0 2 0 3 3
3 3 0 3
23 3 0 3 0 1 3 3 1 0 1 2 1 1 1 1 1 2 0 2 3 3 0 3
5 3 0 2 3 0
3 3 1 1
4 3 0 3 3
7 3 0 3 3 3 0 3
13 3 1 3 0 1 0 1 1 0 1 1 0 2
3 3 0 3
10 3 1 2 0 2 1 3 3 2 3
20 3 1 3 1 3 3 3 3 3 2 0 3 0 1 1 1 2 3 0 2
3 3 0 3
15 3 3 0 2 3 2 0 2 0 3 0 1 3 3 0
3 3 3 0
7 3 0 3 1 0 1 0
25 3 0 3 3 1 3 3 1 1 3 0 3 0 1 3 3 0 3 0 3 0 3 1 2 3
10 3 3 1 1 3 3 3 1 3 3
6 3 0 3 1 2 3
4 3 3 3 2
6 3 1 1 3 0 0
13 3 1 3 0 2 3 2 0 2 0 1 3 3
2 3 3
9 3 0 3 1 3 0 3 0 2
14 3 0 3 0 3 1 0 2 0 0 2 1 2 3
10 3 0 3 3 1 3 0 2 3 0
5 3 1 3 0 0
3 3 3 0
13 3 1 3 1 0 1 3 0 1 2 1 1 0
4 3 3 2 3
48 3 3 1 1 3 3 0 1 1 2 0 3 0 2 2 2 3 0 1 3 3 0 3 2 0 3 0 3 0 0 3 0 1 3 3 3 0 2 1 3 2 0 1 1 1 1 0 1
2 3 2
4 3 3 1 0
10 3 3 0 3 0 3 0 1 2 3
22 3 3 1 3 3 0 1 0 1 3 0 1 2 0 3 1 2 3 0 0 1 3
16 3 0 3 1 1 3 3 0 3 0 3 1 3 1 3 0
1 3
1 3
6 3 3 0 2 1 3
13 3 1 3 0 2 1 3 3 1 3 0 0 0
7 3 0 3 0 1 3 3
9 3 1 3 0 2 0 2 3 0
17 3 0 1 1 3 0 1 2 0 2 3 0 1 1 2 2 3
3 3 1 3
5 3 1 1 3 0
4 3 3 0 0
6 3 3 0 0 1 3
5 3 3 2 0 0
5 3 0 2 1 3
8 3 3 0 0 0 3 3 3
3 3 0 3
6 3 0 3 0 1 2
8 3 0 3 1 0 1 0 2
6 3 3 0 1 1 3
1 3
6 3 0 3 1 2 3
2 3 3
9 3 1 2 1 1 1 3 1 3
2 3 3
21 3 1 1 1 3 0 0 1 3 0 2 0 2 3 0 1 1 1 1 3 3
7 3 3 3 0 0 3 3
23 3 3 0 0 0 1 3 3 3 3 0 1 1 3 0 1 0 0 1 3 3 1 3
2 3 3
14 3 0 3 3 0 2 2 0 3 1 3 3 1 3
7 3 0 3 3 0 1 0
16 3 3 1 3 3 1 0 1 3 3 0 3 0 1 0 2
3 3 0 3
4 3 1 3 0
11 3 1 3 0 2 3 1 3 3 3 0
2 3 3
15 3 3 1 3 3 0 3 0 1 2 3 3 1 0 3
11 3 3 0 0 3 3 2 0 1 3 3
2 3 3
4 3 1 3 0
4 3 0 3 3
8 3 0 3 0 1 3 3 3
5 3 3 1 3 3
15 3 3 0 0 0 3 3 3 1 1 3 0 3 1 3
9 3 0 1 2 1 1 1 1 0
13 3 0 3 1 3 3 0 2 0 3 1 0 2
12 3 1 0 3 3 3 1 3 3 1 3 2
4 3 3 1 3
4 3 0 3 3
13 3 0 3 3 1 3 3 0 3 0 1 2 3
4 3 0 2 3
2 3 3
3 3 3 0
8 3 1 3 0 2 0 3 3
3 3 3 0
3 3 1 3
10 3 3 1 1 1 3 1 3 3 0
5 3 3 0 1 0
11 3 1 3 0 0 1 3 0 2 1 2
8 3 0 3 1 3 1 3 0
5 3 1 1 3 3
14 3 2 0 3 0 0 1 1 3 0 0 1 3 0
3 3 1 3
6 3 0 3 1 3 0
7 3 0 3 0 1 3 3
3 3 3 0
4 3 1 3 0
4 3 3 0 1
14 3 0 3 3 0 1 1 1 1 0 1 3 3 3
2 3 3
7 3 0 2 1 1 3 0
7 3 1 3 0 1 2 3
10 3 1 3 0 2 1 1 1 3 0
5 3 3 1 2 3
7 3 0 3 0 3 1 3
3 3 3 0
3 3 0 3
26 3 3 1 2 3 1 3 3 3 1 3 3 0 3 0 1 2 3 1 3 3 0 3 0 1 2
3 3 3 0
8 3 1 3 0 2 1 1 2
18 3 1 3 0 1 1 1 1 1 2 0 2 3 0 0 1 3 0
8 3 3 1 2 3 3 0 0
7 3 0 2 3 3 3 3
6 3 0 1 0 0 1
11 3 0 2 3 1 3 2 0 0 3 0
2 3 3
4 3 1 1 1
26 3 3 1 1 3 2 1 1 1 1 1 0 1 3 3 3 1 2 0 3 0 2 1 1 3 1
4 3 2 0 3
1 3
3 3 3 0
6 3 1 1 3 0 0
2 3 1
2 3 3
4 3 3 2 0
10 3 0 3 1 3 0 1 1 3 1
4 3 0 1 2
7 3 1 3 0 2 0 3
14 3 1 3 0 1 2 1 3 1 1 3 0 2 3
3 3 0 3
2 3 3
6 3 1 3 0 2 1
1 3
5 3 0 3 0 3
3 3 1 3
2 3 3
4 3 0 3 0
16 3 3 0 2 0 3 1 2 0 1 3 0 2 0 3 0
9 3 0 3 3 0 0 1 3 0
9 3 3 0 1 1 1 1 1 3
2 3 3
23 3 0 3 0 2 3 2 0 3 0 2 0 3 0 1 2 0 3 0 1 2 1 3
3 3 3 0
7 3 3 2 3 1 1 1
4 3 0 3 0
7 3 0 3 1 2 3 1
6 3 0 3 0 1 1
13 3 0 2 3 0 2 0 2 1 3 0 1 3
8 3 0 3 3 3 3 1 3
4 3 3 3 2
3 3 0 3
3 3 3 1
5 3 0 3 0 2
3 3 3 0
9 3 0 2 1 1 3 0 0 3
6 3 3 2 0 1 3
6 3 1 3 0 1 0
11 3 3 3 0 1 1 1 0 2 2 1
8 3 0 3 0 2 3 1 3
1 3
2 3 3
13 3 0 3 0 3 1 0 1 3 3 3 0 0
8 3 0 3 1 3 1 1 3
10 3 3 1 3 3 0 3 3 0 0
2 3 3
10 3 1 2 0 2 0 2 3 0 2
5 3 1 1 1 3
7 3 3 1 3 3 0 3
11 3 1 3 0 2 1 1 1 1 1 1
13 3 0 3 0 1 3 3 1 0 1 2 0 3
2 3 0
6 3 1 3 0 2 2
38 3 3 1 3 3 3 0 2 1 2 1 0 3 3 3 1 3 0 0 3 3 3 3 3 0 3 0 1 3 3 0 3 1 2 3 0 0 0
16 3 0 2 3 1 3 3 3 2 1 3 3 0 2 3 2
7 3 3 1 1 1 1 3
11 3 1 2 0 1 1 1 2 0 3 3
8 3 0 3 1 0 1 2 3
5 3 0 3 0 0
11 3 1 3 0 1 1 2 0 3 1 3
2 3 0
22 3 1 1 3 3 2 0 3 0 1 2 0 3 3 0 2 1 2 0 2 0 3
9 3 3 1 3 3 0 1 3 2
8 3 0 3 3 0 0 1 3
45 3 0 3 0 0 2 3 0 0 3 3 0 1 3 3 0 3 1 3 3 0 0 3 3 0 3 0 1 3 3 0 0 2 0 3 1 0 2 1 3 3 3 3 0 3
7 3 3 1 3 3 0 3
7 3 1 3 1 3 1 3
15 3 3 1 0 0 1 3 3 3 3 1 3 3 0 3
2 3 3
7 3 0 3 1 2 2 3
1 3
4 3 0 3 0
3 3 1 3
6 3 3 0 1 2 3
12 3 0 3 1 2 1 0 1 2 3 0 0
2 3 3
12 3 0 3 0 3 0 3 1 2 1 1 3
8 3 3 1 3 3 0 3 0
7 3 0 1 3 3 3 0
3 3 3 2
7 3 3 1 3 3 3 0
11 3 1 1 1 3 0 1 0 2 3 3
8 3 3 0 1 2 0 3 3
10 3 3 1 3 3 0 3 1 3 0
8 3 0 3 1 2 1 1 1
5 3 0 2 3 0
11 3 1 3 1 0 0 0 0 1 3 0
5 3 0 0 2 3
7 3 1 0 3 3 0 3
2 3 3
2 3 0
8 3 3 1 3 1 3 3 3
3 3 3 0
3 3 3 0
4 3 3 0 0
8 3 1 3 1 3 3 0 1
3 3 0 2
2 3 3
2 3 3
2 3 3
4 3 3 1 3
3 3 1 3
11 3 3 0 0 0 3 3 3 0 0 2
2 3 3
7 3 1 1 3 0 2 0
8 3 1 1 3 3 1 1 3
4 3 1 3 0
5 3 3 1 3 3
2 3 3
10 3 2 0 3 0 2 2 0 3 0
3 3 0 3
4 3 3 3 0
1 3
7 3 1 3 1 3 3 3
3 3 1 3
3 3 3 0
3 3 1 2
8 3 3 0 1 2 3 1 1
9 3 1 3 1 3 3 0 3 0
2 3 3
7 3 3 1 3 3 0 3
3 3 3 0
19 3 0 3 3 2 0 2 0 3 1 2 0 3 1 3 2 0 3 0
7 3 3 0 1 2 1 3
12 3 2 0 3 0 2 0 3 3 1 0 2
7 3 1 0 0 3 0 0
1 3
4 3 0 1 2
4 3 3 1 0
3 3 0 3
7 3 1 3 1 1 2 1
3 3 1 3
3 3 1 3
1 3
24 3 1 2 0 1 1 1 3 0 1 3 3 3 1 0 3 2 2 0 3 1 3 0 2
2 3 3
2 3 3
9 3 0 2 0 1 3 3 0 3
8 3 2 0 1 3 0 1 3
16 3 1 3 1 0 1 1 1 3 3 3 0 2 0 1 3
7 3 3 0 2 1 1 3
9 3 0 2 3 0 1 2 3 2
10 3 3 1 0 3 1 1 2 0 3
13 3 0 3 1 0 1 3 3 1 0 2 2 3
3 3 0 3
5 3 1 3 0 2
2 3 3
20 3 0 3 0 1 3 3 1 0 1 3 3 3 3 1 3 3 1 2 3
9 3 3 0 2 0 0 2 1 0
12 3 0 3 1 1 3 0 1 0 1 3 3
1 3
5 3 0 3 3 3
13 3 0 3 0 3 3 3 0 3 3 1 3 0
16 3 1 3 0 1 1 2 3 0 1 3 3 0 2 3 0
1 3
11 3 0 3 0 1 2 1 2 0 3 0
28 3 0 3 0 2 1 1 3 1 3 0 1 1 1 2 3 2 3 0 0 1 1 3 0 0 1 3 0
7 3 0 2 1 3 0 0
3 3 3 0
5 3 0 3 0 2
8 3 0 3 3 0 1 1 0
4 3 1 3 0
2 3 0
14 3 0 3 1 3 3 1 1 0 0 2 3 0 0
3 3 1 3
12 3 0 3 0 2 0 3 1 1 1 1 0
10 3 3 0 0 0 1 1 2 1 0
29 3 3 1 3 3 3 1 3 3 3 2 0 3 1 0 1 3 3 1 2 2 0 1 1 3 3 0 1 0
3 3 3 2
3 3 0 3
8 3 3 0 2 1 3 1 3
8 3 0 3 1 2 0 3 0
2 3 3
3 3 1 2
11 3 0 3 1 0 2 3 2 0 1 3
5 3 1 1 3 3
2 3 3
9 3 3 0 1 2 3 3 2 1
3 3 3 0
3 3 0 3
12 3 3 0 1 2 3 0 1 2 0 3 0
6 3 0 3 0 1 2
21 3 0 3 3 3 0 3 0 3 0 2 3 0 3 1 0 2 0 2 1 3
12 3 0 3 0 1 3 3 1 1 1 3 3
2 3 3
3 3 0 1
4 3 0 3 0
4 3 3 0 1
5 3 0 3 0 3
4 3 3 0 2
10 3 0 3 0 1 3 3 1 2 3
3 3 3 0
7 3 0 3 1 2 2 3
14 3 1 0 3 3 1 2 0 3 0 2 3 2 3
7 3 1 1 3 1 1 3
8 3 0 1 0 3 2 1 3
14 3 1 3 1 1 2 0 2 3 1 3 3 0 3
19 3 3 1 3 3 0 3 0 3 1 3 0 2 1 3 2 1 3 1
3 3 1 0
8 3 1 3 0 1 2 0 3
2 3 3
7 3 3 1 3 2 1 0
1 3
7 3 3 0 2 1 2 1
2 3 3
2 3 3
2 3 3
15 3 1 1 3 1 1 3 0 2 0 1 0 0 2 0
2 3 3
13 3 3 0 2 1 3 0 1 1 1 2 1 0
6 3 3 1 3 3 3
11 3 1 1 3 0 3 1 2 3 3 0
16 3 0 3 1 0 1 3 2 3 3 3 3 1 2 1 2
9 3 0 3 3 0 0 1 3 3
13 3 0 3 1 2 1 0 1 1 0 3 1 3
19 3 3 1 3 3 0 3 1 3 0 3 1 3 3 0 2 1 3 0
7 3 0 3 1 3 0 1
7 3 3 0 2 2 0 3
2 3 0
1 3
3 3 0 3
4 3 1 3 1
4 3 0 2 3
3 3 1 3
9 3 0 2 1 3 0 1 2 3
2 3 3
23 3 0 3 3 0 0 0 3 3 3 0 2 0 3 0 2 1 1 2 3 0 3 0
9 3 1 0 2 3 0 1 0 0
4 3 3 0 2
1 3
7 3 3 0 0 1 3 0
2 3 3
3 3 3 0
2 3 1
15 3 0 3 3 3 0 3 0 2 3 0 2 3 2 3
6 3 0 3 0 3 0
1 3
25 3 0 3 0 1 3 3 1 0 1 2 1 1 1 2 0 2 3 0 2 2 0 3 0 0
4 3 0 3 0
2 3 0
3 3 0 3
7 3 0 3 0 3 0 3
4 3 0 2 3
9 3 3 0 1 2 0 3 3 2
5 3 0 3 0 2
2 3 2
1 3
29 3 0 3 1 3 0 2 3 0 2 0 1 0 1 3 0 1 2 0 3 0 1 3 3 0 3 3 1 0
4 3 3 0 0
32 3 0 1 3 3 0 3 3 3 3 1 3 3 0 1 2 3 3 1 3 3 1 1 3 0 1 1 1 2 3 1 0
23 3 3 0 0 3 3 0 1 3 3 1 3 0 1 3 3 1 2 3 0 2 0 1
2 3 3
8 3 3 1 3 3 0 0 3
12 3 3 0 1 3 1 1 1 3 3 1 0
17 3 3 1 3 3 3 0 2 0 3 0 1 3 3 3 0 1
7 3 3 1 0 2 3 0
6 3 1 1 3 3 0
3 3 1 3
22 3 0 1 2 3 3 2 0 1 2 1 1 2 0 3 1 2 2 0 2 1 3
10 3 0 3 1 3 1 3 0 2 3
4 3 2 0 3
2 3 3
6 3 0 3 3 3 2
1 3
1 3
22 3 0 1 3 3 3 0 1 3 2 2 0 0 0 1 1 1 1 1 3 1 3
6 3 0 1 0 1 3
13 3 3 1 3 3 3 1 1 1 1 1 2 0
7 3 1 3 0 1 2 3
10 3 3 1 3 3 1 0 2 0 0
4 3 0 2 3
8 3 3 0 1 1 3 2 3
4 3 0 2 3
5 3 1 3 1 3
5 3 3 2 0 0
2 3 3
6 3 0 3 1 2 0
2 3 3
2 3 3
1 3
8 3 1 3 0 3 1 1 1
26 3 3 1 3 3 1 2 1 1 3 0 3 1 2 3 0 0 1 3 0 2 3 2 0 0 3
3 3 3 1
10 3 0 3 0 1 3 2 1 3 3
4 3 2 0 3
9 3 0 2 3 0 1 2 0 3
3 3 3 2
3 3 0 3
14 3 0 3 0 3 3 3 0 1 3 3 1 2 0
2 3 3
8 3 0 1 3 3 1 2 0
3 3 1 0
4 3 1 3 0
2 3 3
4 3 0 2 3
6 3 2 1 0 3 3
13 3 3 1 3 3 1 0 3 1 1 3 1 3
9 3 1 1 3 1 1 1 3 0
1 3
2 3 0
7 3 1 3 0 1 2 3
5 3 3 0 0 3
13 3 3 0 0 1 3 1 3 0 2 2 0 3
3 3 3 0
1 3
3 3 3 0
14 3 3 1 0 3 2 1 1 3 1 3 1 3 3
4 3 3 0 0
7 3 3 2 0 2 0 3
3 3 0 3
3 3 3 0
7 3 0 3 1 2 1 0
7 3 3 0 2 1 3 0
8 3 0 3 1 2 0 3 0
2 3 3
12 3 0 1 2 1 3 0 3 3 0 3 0
3 3 3 0
8 3 0 3 3 3 3 2 1
2 3 3
4 3 1 1 3
4 3 0 3 0
3 3 3 0
2 3 3
1 3
2 3 2
33 3 3 1 3 3 1 2 2 0 3 3 0 3 1 1 1 1 1 1 1 3 3 3 1 1 1 3 3 2 3 1 0 0
2 3 0
2 3 3
4 3 0 3 0
13 3 3 0 1 1 1 1 1 2 1 1 3 0
9 3 0 3 1 2 1 3 3 3
5 3 3 1 3 3
3 3 3 0
23 3 1 1 3 0 1 1 1 1 3 0 1 3 3 1 2 1 1 1 1 2 1 3
4 3 0 3 1
6 3 3 1 2 0 3
4 3 3 0 2
2 3 1
14 3 3 3 3 3 1 2 1 1 3 2 0 2 3
4 3 1 3 0
2 3 3
6 3 0 2 3 1 3
10 3 1 0 0 1 0 2 3 0 3
4 3 1 2 0
4 3 0 3 0
2 3 3
18 3 0 1 2 1 1 3 3 3 3 0 1 2 3 2 0 3 0
5 3 1 1 3 0
7 3 0 3 1 2 3 0
21 3 0 3 0 0 3 0 1 3 3 0 0 1 3 3 0 2 3 0 1 3
12 3 0 3 1 3 1 3 3 1 2 1 0
19 3 0 3 2 0 3 0 2 1 2 0 2 0 3 0 1 3 2 0
11 3 0 3 0 1 3 3 3 3 1 3
12 3 0 1 2 1 3 3 2 0 2 0 3
1 3
22 3 0 3 1 1 3 0 1 3 3 1 0 1 3 3 0 3 1 1 1 1 1
12 3 0 2 0 0 0 0 1 1 2 1 0
5 3 0 3 1 3
5 3 3 0 1 3
3 3 3 0
27 3 0 3 1 0 1 0 1 2 1 2 0 3 0 2 1 1 3 0 0 3 3 3 3 3 1 1
3 3 0 2
2 3 3
2 3 3
7 3 3 1 3 2 0 3
4 3 1 2 0
3 3 3 2
5 3 3 0 2 2
4 3 3 2 0
12 3 0 3 1 0 1 2 1 1 0 1 3
11 3 1 3 0 1 2 0 3 0 2 0
2 3 3
15 3 0 3 1 2 2 0 3 0 1 3 3 3 3 2
3 3 0 1
8 3 0 3 1 3 3 1 3
2 3 3
2 3 0
3 3 3 0
20 3 0 3 1 3 0 3 0 3 3 0 2 1 0 3 0 0 3 2 3
12 3 0 3 0 3 0 1 3 3 3 0 2
8 3 1 0 3 3 1 2 3
3 3 3 2
24 3 3 1 3 3 0 1 3 3 3 1 1 1 1 3 1 2 0 3 1 2 3 3 2
14 3 0 1 2 0 3 1 3 3 1 3 3 3 3
3 3 1 3
11 3 0 3 1 0 1 2 3 0 1 3
3 3 0 1
11 3 0 3 1 2 0 3 0 0 1 3
4 3 0 2 3
3 3 1 3
12 3 0 3 1 2 1 1 1 1 2 3 2
2 3 3
10 3 0 2 2 1 1 1 1 1 0
4 3 1 1 3
4 3 0 3 3
2 3 3
3 3 3 3
5 3 1 3 1 1
6 3 1 3 0 0 0
7 3 0 3 1 2 3 0
3 3 0 3
12 3 1 3 0 2 0 3 0 1 3 3 3
18 3 0 3 0 0 3 0 0 3 0 1 0 3 3 0 3 1 2
23 3 3 1 3 3 3 0 0 0 1 0 1 1 3 2 0 3 0 0 0 1 1 2
8 3 3 3 3 2 0 3 0
7 3 3 3 0 2 0 1
2 3 3
29 3 1 2 0 1 1 3 2 1 2 1 2 1 3 1 3 3 1 2 0 3 0 0 1 3 1 0 1 0
2 3 2
2 3 1
4 3 0 3 0
16 3 3 1 3 3 3 0 1 3 2 3 1 3 2 3 0
2 3 3
8 3 0 3 0 3 0 1 3
8 3 0 3 3 0 1 1 0
4 3 0 3 3
2 3 3
3 3 3 2
6 3 0 3 0 1 2
4 3 3 1 2
3 3 3 0
16 3 0 3 0 3 0 3 1 0 1 0 3 1 3 3 3
8 3 0 3 0 1 3 3 0
5 3 0 2 3 0
7 3 0 2 3 0 1 0
4 3 3 1 3
3 3 3 0
1 3
8 3 3 1 3 3 3 1 1
5 3 0 3 0 2
19 3 3 3 1 3 3 0 3 0 1 3 3 3 0 2 3 1 3 3
20 3 0 2 3 1 3 3 1 3 0 2 0 3 3 3 1 1 3 3 3
4 3 0 2 3
11 3 0 3 1 3 3 1 3 3 3 0
3 3 0 3
1 3
1 3
9 3 3 1 3 3 2 3 0 2
3 3 1 3
3 3 0 3
19 3 3 1 1 1 2 0 3 1 3 3 1 3 3 1 3 3 1 3
4 3 0 3 3
2 3 3
15 3 2 3 1 3 0 3 0 1 1 1 3 0 1 2
12 3 3 0 2 0 3 0 1 3 3 0 3
2 3 0
2 3 3
15 3 0 3 0 1 3 2 3 3 0 1 3 3 1 3
9 3 0 3 0 2 0 3 0 0
26 3 0 3 0 1 1 1 1 1 1 3 2 0 2 0 1 0 0 2 1 3 0 2 1 3 0
5 3 3 1 3 3
4 3 0 2 3
2 3 3
4 3 1 3 1
2 3 3
9 3 0 3 1 2 2 3 1 1
15 3 0 3 0 1 2 1 3 0 0 1 3 3 0 0
11 3 0 3 1 0 1 0 2 1 0 3
9 3 3 0 3 3 0 1 3 3
8 3 0 2 2 0 3 0 2
5 3 0 3 0 3
3 3 3 0
10 3 1 1 2 3 3 0 0 3 0
34 3 0 1 2 1 2 3 1 0 1 2 1 3 0 2 0 0 2 1 1 0 1 3 3 0 3 1 2 1 0 1 3 3 3
7 3 0 3 0 1 0 0
12 3 0 3 0 1 0 2 0 1 3 3 3
3 3 1 3
15 3 2 0 3 0 0 0 1 0 1 3 3 3 3 1
1 3
3 3 3 3
2 3 3
3 3 3 0
9 3 1 3 0 1 1 1 1 0
11 3 0 3 0 1 2 2 0 3 3 0
14 3 3 1 2 1 1 3 2 1 3 2 2 1 3
7 3 3 0 0 3 3 1
1 3
12 3 1 1 3 0 3 0 1 1 1 3 3
5 3 0 3 3 3
2 3 0
10 3 0 3 1 3 2 1 3 0 2
7 3 0 3 1 2 3 0
7 3 0 3 1 2 0 3
3 3 3 2
10 3 1 0 3 3 3 1 3 3 3
2 3 3
3 3 0 3
3 3 3 2
13 3 0 3 3 0 2 0 3 3 1 3 3 0
13 3 3 0 2 0 3 3 1 1 0 2 3 1
10 3 0 3 3 2 3 2 0 3 0
5 3 3 1 3 3
15 3 2 0 3 0 2 3 1 2 1 1 1 1 1 3
5 3 0 3 0 2
3 3 0 3
8 3 3 3 3 3 3 3 3
5 3 0 2 1 3
5 3 0 3 0 2
1 3
4 3 2 0 3
1 3
9 3 0 3 1 3 0 3 1 2
3 3 3 0
1 3
9 3 3 0 2 0 3 1 2 3
2 3 0
1 3
4 3 3 1 2
2 3 3
2 3 3
7 3 0 3 0 1 3 3
2 3 3
7 3 0 3 1 3 3 0
14 3 0 3 0 2 3 0 3 1 0 2 0 0 2
1 3
9 3 1 3 0 1 2 3 0 2
5 3 3 1 3 3
13 3 3 3 1 3 3 1 2 3 0 2 1 2
4 3 1 1 1
29 3 3 3 3 0 1 3 3 3 1 3 3 3 1 3 3 0 1 3 3 0 3 0 1 3 3 1 1 3
15 3 1 1 1 1 1 1 3 1 3 0 2 2 0 3
11 3 0 1 1 3 3 3 1 1 3 0
15 3 2 0 3 0 0 0 2 2 0 3 0 1 3 1
1 3
5 3 0 3 0 3
7 3 1 0 0 2 1 1
8 3 2 0 3 0 0 1 0
2 3 0
3 3 0 1
5 3 0 2 3 0
14 3 0 2 3 2 0 3 0 0 1 3 0 0 3
2 3 3
5 3 3 2 3 3
5 3 1 0 3 3
9 3 3 1 3 3 0 0 2 3
14 3 0 3 0 1 3 3 1 2 1 1 2 0 3
1 3
2 3 3
3 3 0 3
26 3 0 3 0 2 3 0 3 1 3 0 3 0 3 0 2 3 0 3 0 1 1 0 3 1 2
1 3
17 3 0 3 0 1 0 1 3 3 0 3 1 2 2 0 1 0
2 3 0
3 3 0 3
8 3 1 1 3 0 2 3 3
3 3 3 3
15 3 0 3 0 1 1 1 1 1 3 1 1 3 0 2
2 3 3
3 3 0 3
18 3 0 1 2 0 1 3 3 3 1 3 0 3 1 3 0 1 1
4 3 0 2 3
5 3 1 3 0 0
18 3 3 3 1 3 3 0 2 3 1 0 3 1 3 0 0 3 3
2 3 3
6 3 1 3 0 2 0
9 3 3 0 1 1 1 1 0 1
5 3 3 0 0 0
14 3 0 3 0 1 3 3 1 3 1 1 3 1 0
3 3 3 0
1 3
3 3 0 3
14 3 0 3 1 2 3 2 2 0 0 3 0 1 3
9 3 0 3 1 3 0 1 1 1
7 3 2 3 1 3 0 2
3 3 0 3
4 3 0 3 3
5 3 3 0 2 3
5 3 0 2 1 3
3 3 0 3
4 3 0 0 1
16 3 1 1 1 1 2 0 3 3 1 3 3 1 2 3 0
3 3 3 3
11 3 0 3 1 2 3 1 3 3 0 0
13 3 3 2 0 2 1 1 3 3 0 1 1 1
1 3
2 3 1
1 3
14 3 1 3 1 3 3 0 3 0 3 0 1 3 3
5 3 0 3 1 0
10 3 0 3 1 2 2 3 1 2 1
2 3 3
17 3 1 1 3 0 2 0 1 3 3 0 3 3 0 0 1 3
15 3 3 0 0 1 3 0 1 1 0 1 2 1 3 0
5 3 3 2 0 2
5 3 0 3 1 2
1 3
3 3 3 2
7 3 3 1 2 3 0 0
3 3 3 1
3 3 0 3
12 3 1 1 3 0 2 1 1 3 1 3 0
11 3 3 1 3 3 0 1 2 0 1 3
1 3
2 3 3
25 3 0 3 0 3 0 1 1 0 1 3 0 1 1 3 0 3 1 2 1 1 0 0 3 1
5 3 3 2 0 2
32 3 0 1 3 3 1 1 3 1 3 0 2 0 1 2 3 3 1 3 0 2 0 1 1 2 0 3 0 2 2 0 3
6 3 3 1 3 3 3
21 3 1 1 3 3 3 0 2 0 3 0 2 1 1 0 1 3 3 1 3 0
16 3 0 3 1 3 0 1 2 0 3 0 3 1 3 0 2
2 3 3
1 3
20 3 3 1 2 1 3 0 3 0 0 3 0 2 1 2 0 2 3 1 2
5 3 2 0 3 0
6 3 1 1 3 0 1
4 3 3 1 3
4 3 0 2 3
8 3 0 3 1 3 3 0 0
6 3 0 3 0 2 0
3 3 1 2
11 3 0 3 0 3 1 0 2 0 0 2
3 3 3 0
6 3 3 1 2 3 3
4 3 0 2 3
3 3 0 3
7 3 0 3 1 2 0 3
4 3 3 0 0
8 3 3 0 3 3 0 3 3
2 3 3
1 3
3 3 3 0
9 3 0 3 3 0 2 0 3 3
1 3
5 3 0 3 0 3
43 3 3 1 3 3 3 3 1 3 3 3 1 2 3 3 0 3 3 0 3 3 1 3 1 1 1 2 0 2 0 3 1 2 1 1 1 2 0 3 1 2 0 2
10 3 3 0 2 0 1 3 3 3 3
10 3 0 2 3 0 0 3 3 0 3
6 3 1 3 0 1 0
5 3 0 3 0 1
12 3 0 3 0 3 0 1 1 1 1 1 1
2 3 3
2 3 3
6 3 1 1 3 3 3
3 3 3 2
20 3 3 0 1 1 1 2 0 3 1 2 1 3 2 0 3 0 0 1 3
11 3 1 2 0 2 1 3 0 1 1 2
7 3 3 1 2 3 0 0
9 3 0 3 0 3 3 3 1 3
24 3 2 0 3 1 3 3 0 2 3 1 1 3 3 3 1 0 1 1 3 2 2 1 3
3 3 1 3
10 3 0 3 0 1 3 3 1 2 3
2 3 0
4 3 0 3 3
1 3
2 3 3
2 3 3
4 3 3 0 0
8 3 0 1 0 3 1 3 0
8 3 0 3 0 2 3 1 0
9 3 1 3 0 1 3 3 3 1
3 3 0 3
2 3 2
4 3 0 3 3
9 3 3 3 2 0 2 1 3 0
1 3
1 3
4 3 0 1 0
20 3 0 2 3 1 2 3 3 1 3 3 0 1 0 1 0 1 2 1 3
7 3 0 3 1 2 0 3
2 3 3
13 3 0 3 0 3 0 3 3 0 0 1 1 3
2 3 3
15 3 0 3 0 1 3 3 0 1 1 3 3 0 2 3
6 3 0 3 0 1 3
15 3 3 1 3 3 0 0 3 0 1 1 3 2 0 3
1 3
4 3 3 2 3
8 3 3 0 0 3 3 0 3
3 3 3 2
2 3 3
1 3
2 3 3
4 3 3 0 2
11 3 1 1 3 1 3 3 2 0 3 1
10 3 0 3 1 3 1 3 3 1 0
3 3 0 3
2 3 3
4 3 1 1 3
8 3 0 3 0 1 3 3 2
3 3 3 0
19 3 1 3 0 1 1 1 1 2 3 3 1 3 1 3 0 1 1 3
3 3 1 3
10 3 1 3 0 1 0 1 3 3 0
8 3 3 1 3 3 0 3 3
19 3 0 2 3 0 1 1 1 1 0 2 3 1 3 3 1 2 1 3
5 3 1 2 0 0
2 3 0
3 3 0 3
15 3 0 3 1 0 1 3 3 1 0 1 3 3 0 3
3 3 1 3
15 3 3 2 0 2 0 3 0 3 0 1 1 0 0 1
3 3 1 3
4 3 1 1 3
3 3 3 3
17 3 0 2 3 1 2 3 3 0 3 3 1 0 1 3 3 3
4 3 0 3 0
5 3 0 2 3 0
12 3 3 1 0 1 3 3 1 1 1 1 1
3 3 3 2
9 3 3 0 0 0 1 0 0 3
3 3 0 3
4 3 2 0 3
5 3 3 0 3 3
4 3 1 3 0
4 3 0 3 3
13 3 0 0 3 0 1 3 3 3 0 1 2 3
7 3 0 1 0 1 3 0
3 3 3 1
27 3 1 3 0 1 3 0 2 3 2 3 1 3 3 0 3 0 2 2 2 3 0 1 2 1 3 0
3 3 0 3
12 3 3 0 1 2 0 3 3 1 3 3 3
10 3 3 0 1 0 1 1 0 1 0
8 3 0 2 3 1 1 1 3
3 3 1 3
4 3 0 3 3
1 3
2 3 0
8 3 0 3 0 2 0 0 3
1 3
10 3 3 1 1 1 1 1 1 1 3
6 3 1 1 3 3 0
3 3 0 3
3 3 0 3
5 3 0 3 0 2
8 3 0 3 1 3 0 1 1
3 3 1 2
10 3 3 1 3 3 3 1 3 3 0
4 3 1 3 0
4 3 2 0 3
13 3 1 2 1 3 3 0 2 0 0 2 0 3
8 3 2 0 3 3 1 3 0
2 3 3
8 3 3 0 2 0 3 0 3
8 3 0 3 3 3 0 0 3
3 3 0 3
6 3 0 2 3 3 0
5 3 3 0 1 3
3 3 0 3
8 3 3 1 3 1 3 3 3
15 3 3 1 1 1 1 1 1 1 1 1 1 3 1 3
20 3 3 3 0 1 1 2 1 2 3 2 0 0 0 1 1 2 3 0 1
2 3 0
3 3 1 1
4 3 1 2 0
3 3 1 3
10 3 0 3 0 1 1 1 1 1 1
3 3 1 3
3 3 1 2
15 3 0 3 1 3 3 1 3 3 0 3 0 1 3 3
8 3 1 3 1 3 3 0 3
4 3 1 1 1
3 3 3 0
6 3 0 1 2 2 3
4 3 3 0 0
2 3 3
4 3 0 3 0
3 3 0 3
3 3 3 2
1 3
1 3
25 3 3 1 3 3 3 1 0 1 3 3 0 3 0 1 2 0 2 0 1 3 3 3 2 0
7 3 0 3 0 1 3 2
1 3
7 3 3 1 3 3 3 0
36 3 0 3 0 1 2 3 1 3 0 2 2 3 1 2 2 3 1 3 3 1 2 3 0 2 0 1 2 1 1 1 1 1 1 2 3
3 3 1 3
2 3 3
8 3 3 3 0 3 3 1 3
3 3 1 3
9 3 0 3 0 3 0 1 3 3
5 3 2 3 0 1
2 3 3
30 3 0 3 0 1 3 3 3 3 1 3 3 3 0 2 0 1 2 3 0 3 0 1 3 3 1 1 1 1 3
4 3 1 3 0
1 3
8 3 2 0 3 0 2 0 3
3 3 1 3
1 3
4 3 3 0 1
2 3 3
17 3 3 1 3 3 1 2 2 3 2 3 1 1 3 3 1 3
10 3 3 0 0 1 3 0 1 2 0
2 3 3
3 3 3 0
20 3 3 0 0 3 0 0 1 2 3 0 1 3 1 1 3 0 1 1 2
3 3 0 3
3 3 3 0
8 3 0 3 1 2 1 3 2
1 3
4 3 0 3 3
10 3 1 1 3 3 1 3 1 2 3
5 3 3 1 0 3
10 3 3 1 3 0 0 3 0 0 2
4 3 2 0 3
3 3 1 3
8 3 0 3 3 0 0 1 3
5 3 0 2 3 0
9 3 0 1 2 0 3 0 3 3
31 3 3 0 2 1 1 1 3 0 3 3 0 2 3 0 1 3 3 3 3 0 3 0 3 1 3 1 1 3 3 1
7 3 0 3 1 2 2 3
2 3 3
6 3 0 3 1 3 0
31 3 3 0 1 2 0 3 0 1 3 1 2 0 3 1 0 1 2 1 2 0 3 0 1 3 3 0 1 3 3 3
12 3 3 1 3 3 1 3 3 2 0 0 0
3 3 3 2
3 3 3 2
2 3 3
3 3 0 3
5 3 1 1 3 3
2 3 3
2 3 0
3 3 0 3
5 3 0 2 3 0
2 3 3
4 3 1 3 0
5 3 0 2 3 0
10 3 1 3 1 3 1 3 3 1 3
2 3 3
6 3 3 0 0 1 3
16 3 0 2 3 0 1 1 1 1 1 1 0 1 1 0 3
8 3 3 0 0 1 3 0 2
6 3 0 3 1 3 3
3 3 1 3
3 3 0 3
25 3 3 0 2 0 3 1 0 2 1 2 1 1 1 3 0 0 1 3 1 3 3 0 2 3
12 3 3 1 0 2 2 3 0 3 1 3 3
8 3 0 1 2 2 0 3 0
10 3 3 1 3 3 3 1 3 3 3
5 3 0 3 0 2
4 3 0 3 3
4 3 3 3 2
13 3 0 2 3 0 1 2 0 3 0 3 3 1
4 3 0 2 3
4 3 0 1 2
2 3 3
30 3 0 3 1 2 2 0 3 0 3 0 1 3 3 0 2 1 0 1 3 3 0 3 3 0 1 2 3 2 3
4 3 0 3 3
5 3 3 3 1 3
15 3 1 3 1 3 1 1 1 1 2 0 2 3 0 0
5 3 1 1 3 0
12 3 0 2 3 0 2 1 1 3 1 0 3
12 3 0 3 1 2 2 0 1 2 2 1 3
17 3 0 2 3 1 1 3 0 1 1 1 0 1 3 3 3 3
10 3 0 1 3 3 1 2 0 3 0
14 3 0 3 0 3 0 1 2 0 3 0 2 3 3
6 3 0 3 0 2 3
1 3
13 3 0 1 3 3 3 2 1 3 3 0 3 3
4 3 0 2 3
3 3 0 1
14 3 1 3 0 1 3 0 0 1 3 0 2 3 2
2 3 3
4 3 0 3 0
9 3 3 1 3 3 0 1 3 3
6 3 3 1 0 0 1
13 3 3 1 3 3 3 1 0 2 1 1 0 0
9 3 0 3 0 2 3 1 1 2
4 3 0 3 3
4 3 0 3 3
25 3 3 1 3 3 1 3 0 2 1 3 1 3 3 0 2 3 3 0 1 1 1 1 1 0
8 3 0 3 0 3 2 0 2
4 3 0 2 3
11 3 0 3 1 0 1 3 3 0 3 3
3 3 1 3
1 3
13 3 1 3 3 0 1 3 3 3 2 3 1 1
3 3 0 3
4 3 3 2 1
2 3 3
3 3 1 3
25 3 0 3 0 2 3 1 3 3 0 1 2 3 0 1 3 3 0 2 3 0 2 2 0 3
8 3 0 3 0 2 1 2 3
5 3 3 0 0 0
1 3
4 3 1 0 0
2 3 3
6 3 3 2 0 2 3
3 3 1 2
2 3 3
11 3 0 3 0 1 3 1 3 0 2 0
2 3 3
2 3 3
5 3 0 2 1 3
2 3 3
2 3 3
17 3 0 3 0 0 3 1 2 1 0 3 3 1 3 0 3 2
3 3 1 3
4 3 0 3 0
4 3 0 3 0
9 3 3 0 2 2 0 3 0 2
3 3 0 3
4 3 0 3 1
6 3 0 1 1 1 0
6 3 0 3 0 2 3
12 3 1 3 1 3 0 0 1 3 3 0 3
7 3 3 0 0 1 1 3
7 3 2 0 3 3 1 3
9 3 3 2 0 2 2 3 1 3
2 3 1
1 3
2 3 3
9 3 1 3 0 2 1 1 1 3
12 3 1 1 1 3 0 2 0 2 1 3 0
6 3 3 0 1 2 3
2 3 3
10 3 3 0 2 0 3 1 3 0 3
4 3 1 3 1
8 3 3 0 0 3 3 0 3
2 3 3
12 3 3 0 2 0 0 0 1 2 0 1 3
16 3 0 3 1 3 3 1 0 2 3 0 1 0 2 3 2
2 3 0
2 3 0
2 3 3
10 3 3 0 2 2 0 3 1 0 3
10 3 1 3 1 3 3 1 3 1 3
21 3 0 3 3 3 1 0 3 3 3 3 0 1 3 3 0 3 0 3 1 3
6 3 0 3 0 2 3
7 3 3 0 2 1 3 0
9 3 3 0 2 2 0 0 3 1
25 3 0 3 0 3 3 1 3 3 0 2 3 0 2 3 1 3 3 0 3 0 1 2 0 3
3 3 0 3
6 3 3 2 0 0 2
2 3 3
5 3 0 2 1 3
15 3 0 3 1 0 2 0 0 2 0 3 1 3 1 3
7 3 2 0 3 0 0 3
7 3 1 3 0 3 3 1
5 3 0 3 1 3
6 3 0 3 1 2 3
6 3 3 1 3 3 3
3 3 3 0
3 3 0 3
2 3 3
1 3
8 3 0 3 0 3 0 2 0
2 3 3
32 3 1 1 3 1 3 1 3 3 3 0 2 0 1 2 3 3 0 0 0 0 0 3 0 1 2 0 3 0 0 1 3
9 3 0 0 3 1 2 1 1 0
14 3 1 1 3 1 2 3 3 2 0 0 1 3 0
8 3 3 0 0 1 3 1 0
11 3 3 1 3 3 0 2 3 1 3 3
13 3 0 3 1 0 1 3 3 0 3 1 0 1
1 3
5 3 3 0 2 3
13 3 1 3 1 1 3 1 3 0 2 1 1 1
10 3 0 3 1 0 1 2 3 3 0
2 3 3
7 3 1 0 3 3 0 2
2 3 3
13 3 1 1 1 1 3 0 3 0 3 2 1 2
4 3 1 3 1
6 3 1 3 0 1 1
9 3 3 0 0 0 3 0 2 3
7 3 0 3 0 2 3 3
10 3 0 3 0 1 3 3 0 2 3
4 3 0 2 3
20 3 3 1 1 2 0 3 1 2 1 3 1 1 1 1 1 3 3 2 1
2 3 0
4 3 1 3 0
4 3 2 0 3
7 3 0 0 2 3 0 2
20 3 0 3 1 2 0 1 3 0 1 0 1 1 0 3 1 3 3 0 3
3 3 1 2
23 3 0 3 1 2 1 1 1 1 1 3 2 2 0 3 3 1 3 3 3 0 2 3
9 3 0 2 3 1 3 3 3 1
16 3 1 1 3 0 3 0 3 0 2 0 0 1 0 1 0
4 3 0 2 3
13 3 3 1 3 3 3 0 1 3 0 1 3 3
2 3 3
6 3 0 1 0 1 3
10 3 1 3 1 3 1 3 1 1 1
6 3 0 3 0 0 3
4 3 0 2 3
16 3 0 3 2 0 3 1 3 3 0 3 0 1 3 3 3
2 3 3
3 3 0 3
6 3 2 0 1 1 3
16 3 0 1 2 2 3 1 2 1 1 1 2 0 3 0 1
3 3 3 0
17 3 0 3 1 0 2 3 1 3 3 3 1 3 3 1 3 0
14 3 0 3 1 2 1 3 0 1 3 3 0 3 0
4 3 3 0 2
3 3 0 3
2 3 3
4 3 1 1 3
12 3 3 0 2 1 1 3 0 3 0 0 1
7 3 3 1 2 3 0 3
4 3 1 1 3
16 3 0 3 1 0 2 2 2 3 0 2 0 3 1 2 3
9 3 0 3 0 1 3 3 3 0
25 3 3 3 3 3 1 3 3 0 3 1 1 3 3 1 0 1 3 3 0 3 0 2 0 3
8 3 0 3 3 3 3 3 1
8 3 3 0 0 0 3 3 3
3 3 0 3
1 3
12 3 0 3 1 0 2 3 3 3 0 1 1
23 3 3 0 2 0 3 3 1 2 1 1 0 2 0 2 1 0 1 2 1 3 3 3
2 3 3
1 3
8 3 3 1 1 3 1 3 0
13 3 3 1 1 1 3 0 3 0 1 0 3 1
12 3 0 3 0 3 0 1 1 3 2 0 3
9 3 0 3 3 0 2 1 1 3
19 3 1 3 1 1 1 1 2 1 3 0 0 0 3 3 3 0 2 3
10 3 0 3 0 1 2 0 3 0 2
20 3 0 3 0 1 2 1 1 1 2 0 3 3 0 1 3 0 1 2 3
1 3
8 3 1 1 1 1 1 2 3
14 3 0 2 3 0 0 0 1 3 3 3 3 0 2
3 3 1 3
27 3 0 3 1 3 0 2 0 3 3 0 0 1 3 1 3 3 3 1 2 1 3 1 1 1 3 0
2 3 3
4 3 1 3 0
4 3 1 1 3
3 3 0 3
2 3 3
2 3 3
5 3 3 0 2 3
2 3 3
14 3 0 3 1 0 1 2 2 0 3 3 3 1 2
19 3 0 3 0 1 3 3 1 1 3 0 2 3 0 2 0 3 0 3
5 3 0 3 0 3
5 3 3 3 3 3
10 3 3 1 0 2 1 3 0 3 3
3 3 1 3
8 3 3 0 0 1 3 0 2
7 3 3 1 3 3 0 3
5 3 3 2 0 0
13 3 0 3 1 0 1 2 3 3 1 3 2 3
11 3 0 3 0 1 2 3 1 0 3 3
7 3 1 2 0 0 1 3
12 3 3 1 0 0 2 0 3 1 3 0 3
12 3 0 3 1 2 1 2 0 3 1 2 1
12 3 0 3 0 1 2 1 2 3 1 2 2
8 3 3 2 3 1 0 1 3
2 3 3
2 3 0
6 3 0 3 0 3 0
7 3 3 0 0 1 3 0
6 3 1 0 3 3 3
4 3 0 3 3
7 3 3 0 1 2 0 3
3 3 0 2
33 3 3 2 0 0 1 1 3 3 0 1 2 3 0 0 1 3 1 3 3 3 1 3 3 0 1 2 0 2 3 2 0 3
3 3 3 0
2 3 1
5 3 3 1 3 3
2 3 0
19 3 3 0 2 0 3 1 2 1 0 0 1 1 1 3 1 1 0 1
12 3 3 1 3 0 3 1 2 1 3 0 1
2 3 3
10 3 0 3 3 3 3 0 1 1 1
13 3 0 3 0 1 3 0 3 3 3 3 2 1
3 3 3 0
7 3 3 1 3 3 3 2
2 3 3
2 3 3
14 3 1 0 2 1 1 0 1 3 3 0 1 3 3
8 3 0 2 3 0 2 0 3
4 3 1 1 1
4 3 3 2 0
3 3 0 3
8 3 1 3 0 2 2 0 3
3 3 0 3
11 3 3 2 3 2 0 3 0 0 1 3
8 3 0 2 3 0 1 1 0
4 3 0 3 0
1 3
21 3 3 0 1 0 0 1 3 3 1 3 3 0 1 1 1 1 1 2 0 3
6 3 1 1 3 0 3
2 3 3
5 3 0 3 0 3
3 3 3 0
11 3 1 3 0 2 0 3 0 1 0 3
6 3 0 3 0 2 1
4 3 3 3 2
4 3 0 2 3
11 3 2 3 0 1 3 3 1 3 3 0
3 3 1 3
4 3 1 3 0
6 3 0 1 2 2 0
11 3 0 3 0 3 1 3 3 1 0 3
20 3 3 1 3 3 0 3 0 1 2 1 1 1 1 1 2 3 2 0 0
4 3 1 3 0
6 3 0 3 0 1 3
5 3 1 1 1 1
2 3 0
7 3 2 0 1 3 0 0
6 3 3 0 0 1 3
2 3 3
3 3 0 3
5 3 0 1 3 3
3 3 0 3
5 3 1 3 1 3
2 3 3
5 3 3 0 1 3
3 3 3 0
3 3 0 3
1 3
1 3
3 3 3 0
10 3 3 1 2 3 0 1 0 1 3
14 3 3 1 3 3 0 3 3 0 2 1 3 0 2
6 3 0 3 0 3 0
5 3 0 3 0 3
19 3 3 2 1 1 2 2 0 2 2 1 1 3 1 3 3 3 0 3
5 3 0 3 3 3
44 3 1 3 1 3 3 2 0 3 0 1 2 1 3 0 0 0 3 1 3 0 1 3 3 0 3 0 1 3 3 0 3 1 2 0 1 0 1 3 3 0 2 3 0
3 3 0 3
6 3 0 2 3 0 0
3 3 0 3
2 3 2
20 3 1 3 1 3 3 3 0 0 1 3 0 0 3 3 1 1 3 3 3
16 3 0 3 1 2 2 1 2 1 2 0 3 1 1 1 3
6 3 0 3 0 3 0
1 3
10 3 0 3 0 3 0 0 3 1 0
3 3 3 1
6 3 3 0 0 3 3
5 3 3 0 2 2
12 3 3 0 1 1 3 3 2 2 1 1 3
8 3 0 3 0 3 1 1 3
9 3 0 3 0 1 0 1 3 3
1 3
19 3 0 3 1 0 1 2 2 0 3 0 3 0 1 1 3 0 3 0
7 3 3 0 2 0 2 3
5 3 3 0 1 3
1 3
2 3 3
5 3 1 3 3 0
6 3 0 3 1 2 3
3 3 1 3
8 3 0 3 0 3 0 1 2
2 3 3
15 3 3 1 0 0 1 3 3 3 2 0 3 0 0 0
2 3 3
3 3 3 3
6 3 1 3 0 1 0
4 3 1 2 3
3 3 0 3
5 3 0 3 1 3
6 3 1 1 3 0 0
3 3 3 2
4 3 0 3 0
3 3 3 0
5 3 0 3 0 3
18 3 1 1 3 0 2 0 3 3 2 1 3 3 0 1 0 0 1
4 3 2 0 3
6 3 0 3 0 3 1
4 3 0 1 0
4 3 0 3 0
16 3 3 1 3 3 3 1 2 3 3 3 0 0 1 3 0
5 3 0 3 3 0
3 3 1 3
3 3 0 2
4 3 1 1 1
12 3 3 2 3 1 3 1 3 0 0 1 3
3 3 3 0
4 3 0 3 0
4 3 3 0 2
11 3 1 3 0 2 1 2 0 2 1 2
2 3 3
6 3 3 1 3 3 3
9 3 0 3 1 2 0 3 0 0
4 3 0 2 3
7 3 0 3 1 2 1 3
10 3 0 3 0 3 3 0 0 1 3
5 3 3 0 1 1
2 3 3
33 3 3 2 0 2 3 1 3 3 0 3 0 3 0 3 1 2 1 1 2 3 1 3 3 3 0 2 0 1 3 3 0 2
1 3
9 3 0 3 0 1 3 3 0 2
20 3 2 0 3 0 1 2 3 0 1 3 1 1 0 1 2 1 1 1 1
16 3 0 1 2 3 0 1 2 3 2 3 0 3 1 2 1
4 3 0 3 3
16 3 3 0 3 1 2 0 0 0 2 2 0 3 0 0 0
3 3 3 2
11 3 0 2 3 0 2 0 3 0 0 3
3 3 1 3
5 3 0 3 1 3
1 3
10 3 1 1 0 3 1 1 2 0 3
7 3 0 2 0 0 0 0
10 3 0 3 1 2 1 1 1 3 1
5 3 1 3 0 1
21 3 3 1 3 3 0 3 1 2 1 1 0 1 1 1 2 2 0 3 1 3
1 3
5 3 0 3 1 3
8 3 1 3 0 0 0 1 1
2 3 3
5 3 0 3 1 3
10 3 3 0 2 0 2 3 2 0 3
8 3 0 2 1 1 1 3 0
4 3 0 3 0
6 3 3 1 3 3 3
1 3
3 3 1 3
8 3 0 3 1 3 3 2 0
14 3 0 3 3 0 0 1 3 0 1 1 2 0 3
22 3 3 1 3 3 3 2 0 1 2 0 0 1 1 2 0 3 3 0 2 3 0
10 3 0 3 3 3 0 3 0 2 3
17 3 3 1 3 3 0 1 3 3 1 1 3 3 0 0 1 3
11 3 0 2 1 3 1 3 3 1 0 0
11 3 0 2 1 3 1 3 3 0 1 2
11 3 1 1 3 0 1 0 1 3 3 3
12 3 3 0 1 2 0 3 0 2 1 1 3
6 3 0 3 1 0 2
1 3
18 3 1 1 3 3 1 3 3 0 3 1 3 3 1 3 2 0 3
16 3 3 0 0 1 3 0 1 1 1 2 3 1 3 1 0
4 3 0 3 3
7 3 3 0 0 0 1 0
9 3 3 0 2 0 3 0 3 3
3 3 1 3
7 3 3 1 3 3 1 3
4 3 1 3 0
12 3 3 1 3 3 3 0 0 0 3 3 3
4 3 0 3 0
10 3 0 3 0 2 1 1 2 1 0
3 3 0 3
16 3 0 1 1 3 2 1 1 2 0 3 0 3 0 2 1
11 3 1 3 1 0 3 3 3 0 2 3
3 3 3 0
3 3 2 0
9 3 0 3 3 2 0 1 0 3
5 3 1 3 0 2
1 3
6 3 1 3 0 2 0
10 3 0 3 0 3 0 3 1 2 3
2 3 3
3 3 0 3
3 3 2 3
4 3 3 0 2
4 3 1 3 0
14 3 0 3 3 1 0 2 2 0 3 0 2 3 2
32 3 0 3 0 2 0 3 0 2 0 3 0 1 2 0 2 0 3 0 3 3 0 1 2 0 3 0 1 1 3 0 3
3 3 1 0
5 3 0 1 2 1
1 3
2 3 3
8 3 1 1 3 0 0 1 3
3 3 3 0
9 3 2 0 3 0 1 2 0 3
15 3 3 1 3 0 1 1 2 1 2 1 3 3 0 3
10 3 0 3 0 3 3 1 3 3 3
1 3
35 3 0 2 3 1 0 2 1 2 2 0 3 0 2 1 3 2 0 1 1 1 2 0 1 2 0 3 1 2 1 1 1 1 0 2
9 3 0 3 1 2 2 0 2 3
3 3 0 3
8 3 1 1 3 1 3 3 3
4 3 0 1 1
5 3 1 1 3 0
3 3 3 0
4 3 3 2 1
3 3 1 3
21 3 1 3 0 2 2 0 3 0 1 1 0 1 3 3 3 3 0 0 1 3
3 3 0 3
14 3 0 3 0 1 3 1 0 1 3 0 1 0 1
1 3
2 3 3
4 3 1 3 1
7 3 0 3 1 2 1 1
4 3 3 0 0
2 3 3
3 3 0 3
3 3 0 3
2 3 3
6 3 1 3 0 1 0
3 3 1 3
2 3 3
3 3 0 3
1 3
11 3 3 1 3 3 1 2 0 2 0 3
17 3 3 1 2 2 0 3 3 0 1 1 3 0 1 0 0 3
6 3 0 3 1 1 3
1 3
4 3 2 0 3
9 3 0 3 0 3 0 1 1 0
6 3 0 3 1 2 1
4 3 1 1 3
2 3 3
13 3 3 1 1 1 2 2 3 1 3 0 3 0
13 3 1 1 3 1 1 3 1 3 3 1 2 3
2 3 1
8 3 3 0 2 1 3 0 0
7 3 0 3 0 2 3 0
1 3
3 3 1 3
2 3 2
3 3 0 3
2 3 0
4 3 3 2 0
1 3
2 3 0
13 3 3 0 1 3 2 0 3 1 2 3 1 0
4 3 1 1 3
4 3 0 3 3
28 3 0 1 2 0 3 0 2 3 0 3 0 1 3 3 1 2 1 2 0 3 1 0 1 2 1 3 0
4 3 0 1 2
12 3 0 3 0 3 0 3 0 3 0 2 0
5 3 3 0 2 0
17 3 0 3 1 0 1 2 2 1 2 1 3 1 3 0 0 3
10 3 0 3 1 1 3 3 1 3 3
4 3 0 3 3
7 3 0 3 1 3 3 2
7 3 3 1 3 3 0 2
3 3 3 2
15 3 3 0 1 1 1 1 1 2 0 2 3 0 0 3
7 3 0 3 0 3 0 2
31 3 3 1 3 3 0 1 2 1 0 1 3 1 3 3 0 1 1 0 2 0 1 2 3 0 2 3 3 1 2 3
10 3 1 3 1 3 3 1 2 3 0
6 3 0 3 1 3 3
2 3 3
6 3 1 1 3 3 3
13 3 0 3 1 0 1 2 1 1 1 1 1 3
3 3 3 0
2 3 3
1 3
1 3
14 3 1 1 1 1 0 3 0 3 1 0 1 3 3
11 3 3 0 0 3 0 0 0 1 1 3
8 3 3 0 2 0 3 0 2
1 3
3 3 1 2
7 3 1 1 3 0 3 0
7 3 0 0 3 1 3 3
2 3 0
6 3 3 1 3 3 3
3 3 0 1
18 3 3 0 2 2 3 0 2 0 3 2 0 3 0 1 2 1 3
1 3
4 3 1 0 0
3 3 0 3
8 3 2 0 1 1 3 3 3
4 3 3 1 0
7 3 0 3 1 3 1 3
5 3 1 3 0 0
2 3 3
7 3 0 2 3 1 3 3
2 3 3
15 3 3 1 3 3 0 2 0 3 1 3 3 2 3 1
5 3 0 2 3 0
11 3 3 0 1 2 0 3 1 3 3 2
8 3 0 3 1 3 1 3 3
4 3 1 3 0
10 3 0 1 0 1 3 3 0 3 3
3 3 3 1
10 3 3 1 1 1 1 1 2 0 3
12 3 0 3 1 0 1 2 2 0 3 0 3
21 3 1 1 1 3 0 0 0 3 3 3 0 3 1 2 3 0 2 0 0 0
5 3 3 1 0 0
6 3 0 3 0 2 1
9 3 0 3 1 2 0 1 1 3
3 3 0 3
8 3 3 1 3 3 0 1 2
3 3 3 0
3 3 1 2
2 3 0
2 3 3
8 3 0 3 0 2 0 1 3
6 3 0 3 1 3 3
13 3 0 1 0 1 2 0 3 1 1 3 2 0
5 3 3 1 0 3
10 3 0 3 0 2 1 0 1 3 3
2 3 3
3 3 1 3
4 3 3 0 2
4 3 3 1 2
11 3 3 0 0 0 0 0 2 2 0 3
4 3 0 3 0
9 3 0 2 3 1 3 0 2 3
4 3 3 0 2
3 3 0 3
8 3 0 3 0 1 2 3 0
10 3 3 1 0 0 2 3 1 1 1
2 3 3
8 3 0 3 3 0 2 0 3
9 3 0 3 0 1 3 0 2 3
8 3 0 3 0 0 0 3 3
9 3 1 3 0 0 3 3 0 3
10 3 3 0 1 1 2 0 1 1 3
3 3 3 3
7 3 0 1 2 3 3 2
5 3 3 1 3 3
10 3 0 3 0 1 3 2 0 0 0
9 3 3 0 1 1 1 2 1 3
7 3 1 1 3 3 3 0
14 3 3 0 0 1 3 0 2 0 3 1 2 1 0
1 3
10 3 0 3 1 3 3 1 1 1 2
5 3 0 2 3 0
5 3 0 2 3 0
3 3 3 2
20 3 1 3 0 3 3 3 2 3 0 3 1 3 1 3 1 3 3 1 3
8 3 3 0 0 0 1 0 3
7 3 3 0 1 2 3 2
4 3 2 0 3
12 3 3 0 2 2 0 2 2 1 2 1 3
14 3 1 3 2 0 1 1 1 2 3 1 2 0 3
3 3 3 0
18 3 0 3 0 1 3 3 0 1 0 1 3 2 3 3 3 3 3
6 3 3 0 1 2 3
3 3 1 3
3 3 1 3
4 3 0 3 0
4 3 0 3 3
5 3 2 0 3 0
2 3 3
2 3 3
2 3 3
27 3 0 3 1 2 1 1 1 2 1 3 0 2 0 1 2 3 0 0 3 0 2 1 2 0 2 3
3 3 3 0
3 3 1 3
9 3 1 3 0 0 1 1 3 0
10 3 1 1 3 0 2 3 1 3 1
3 3 0 3
7 3 0 2 3 0 1 1
2 3 3
3 3 0 1
2 3 0
12 3 3 2 0 2 0 2 3 2 0 0 3
8 3 2 0 3 0 0 1 3
1 3
10 3 3 0 2 1 0 3 3 0 2
5 3 0 3 0 3
7 3 0 0 2 0 1 3
6 3 0 3 1 3 0
43 3 3 0 1 1 1 1 1 3 0 2 3 1 0 3 3 3 0 2 1 0 3 3 1 0 1 3 3 1 2 3 0 0 0 1 3 3 3 0 2 3 0 1
3 3 3 0
5 3 0 2 3 0
4 3 0 3 0
3 3 0 3
7 3 3 0 0 1 3 0
6 3 3 0 2 0 2
1 3
9 3 0 3 0 3 0 1 1 2
2 3 3
2 3 3
2 3 2
6 3 0 3 1 3 3
23 3 0 3 3 1 0 1 3 3 0 0 3 1 0 1 3 3 0 3 0 1 3 2
7 3 0 3 3 2 1 3
6 3 3 0 1 3 0
2 3 3
9 3 0 3 1 2 3 0 0 3
16 3 0 3 1 2 0 3 1 3 3 0 1 2 0 1 3
12 3 3 0 2 2 0 1 1 3 0 1 0
27 3 0 3 3 3 1 2 1 0 1 3 1 3 2 1 3 0 2 3 2 0 1 3 1 3 1 2
7 3 0 3 1 2 1 3
9 3 3 1 3 3 0 1 2 0
3 3 0 3
2 3 1
14 3 0 3 0 3 1 2 1 2 3 1 2 1 3
4 3 1 3 1
2 3 3
3 3 0 3
14 3 0 3 1 3 3 3 3 3 0 0 2 0 3
3 3 1 3
4 3 0 2 3
17 3 3 2 0 1 2 0 3 1 3 3 3 1 3 3 0 3
7 3 0 3 1 2 0 2
11 3 3 0 2 0 3 1 2 3 0 0
2 3 3
19 3 3 0 2 0 3 1 0 1 3 3 0 3 1 3 3 3 0 3
3 3 0 3
10 3 1 1 3 0 3 1 3 3 2
5 3 0 2 3 3
2 3 2
3 3 3 1
3 3 1 3
13 3 1 1 3 3 0 3 0 2 0 0 2 0
1 3
7 3 3 0 1 1 1 0
21 3 0 3 0 3 0 1 0 3 3 3 2 3 0 3 0 1 2 3 0 1
10 3 1 0 3 3 3 2 0 0 0
3 3 3 0
15 3 0 2 1 1 3 3 1 3 0 2 0 1 0 3
7 3 3 0 0 1 3 0
2 3 3
2 3 3
4 3 0 3 3
15 3 3 0 2 0 3 1 2 1 2 3 2 3 1 0
9 3 3 1 2 1 1 2 0 3
3 3 1 3
3 3 3 0
3 3 1 2
16 3 0 2 1 0 2 1 0 1 1 1 1 3 0 1 1
9 3 3 1 3 1 2 0 3 0
7 3 0 3 0 1 3 3
2 3 3
16 3 0 2 3 0 2 1 2 0 2 2 2 1 1 3 1
2 3 3
8 3 3 0 2 0 3 0 3
3 3 0 3
8 3 3 1 1 0 0 3 0
9 3 0 1 3 3 0 2 2 3
3 3 3 0
17 3 0 3 0 1 0 2 3 0 1 3 3 0 3 1 3 3
7 3 1 3 0 0 1 3
2 3 3
9 3 0 2 3 1 1 1 1 1
7 3 0 3 1 2 1 3
2 3 0
9 3 0 1 2 1 1 3 3 0
3 3 0 3
7 3 1 3 0 1 1 3
10 3 0 1 0 3 2 0 3 3 0
3 3 0 3
6 3 1 3 1 3 3
2 3 3
3 3 0 3
4 3 3 1 1
9 3 0 3 1 2 1 1 1 3
3 3 0 3
8 3 0 3 0 3 1 2 3
24 3 1 3 3 2 1 1 1 2 0 3 1 2 3 0 1 2 0 1 3 3 3 2 3
2 3 3
13 3 0 3 1 3 0 3 0 1 0 0 2 1
7 3 3 2 0 2 0 1
22 3 0 3 0 0 3 0 1 3 3 1 3 3 0 2 0 3 1 2 0 3 0
19 3 0 3 0 0 3 1 2 3 0 2 0 1 3 3 0 1 0 0
3 3 0 1
3 3 1 2
16 3 3 1 3 3 1 0 1 2 0 3 1 1 1 1 3
5 3 0 3 1 1
8 3 0 3 0 1 3 1 1
5 3 3 2 0 0
15 3 3 1 3 3 0 1 3 3 1 2 1 1 2 0
1 3
28 3 3 1 3 3 3 1 1 1 1 1 1 0 3 3 1 2 1 1 3 3 3 3 3 0 0 1 3
6 3 1 1 1 3 0
6 3 1 0 1 1 3
1 3
5 3 0 3 1 2
3 3 0 3
8 3 0 0 2 2 1 3 0
3 3 3 0
4 3 1 3 0
6 3 0 3 1 2 3
9 3 2 0 3 1 1 0 3 3
11 3 3 1 3 3 1 2 2 1 3 0
7 3 3 1 3 3 3 0
15 3 0 2 1 1 2 1 2 0 3 1 3 0 2 3
9 3 1 3 0 2 3 1 3 0
7 3 1 1 1 1 2 0
17 3 1 3 3 1 3 0 3 1 3 3 1 3 3 1 0 2
2 3 3
3 3 1 2
8 3 0 3 1 2 1 1 3
8 3 1 3 1 3 3 3 2
3 3 0 3
10 3 0 3 1 2 1 1 2 0 3
12 3 1 1 3 1 1 0 3 2 0 1 3
3 3 3 1
5 3 3 1 2 3
2 3 3
7 3 3 3 1 3 1 3
4 3 1 2 0
7 3 0 3 0 1 3 2
3 3 0 3
22 3 0 3 1 0 2 3 0 3 0 1 3 3 0 0 3 0 1 0 2 2 3
14 3 0 2 3 0 1 1 1 2 3 1 3 3 3
11 3 0 3 3 0 0 3 0 0 1 0
7 3 0 3 1 2 1 0
1 3
3 3 3 0
9 3 3 2 3 1 1 1 1 3
8 3 3 1 3 3 0 3 3
10 3 0 3 0 1 0 1 2 1 3
6 3 0 3 0 1 2
8 3 3 1 3 3 1 3 3
2 3 3
4 3 0 3 0
11 3 0 3 0 1 3 3 0 1 2 0
2 3 0
4 3 0 3 0
2 3 3
4 3 3 3 2
5 3 0 0 0 3
2 3 1
18 3 0 3 3 0 2 3 1 3 0 1 3 3 0 3 1 2 1
9 3 0 3 1 2 1 3 1 0
3 3 0 3
2 3 3
7 3 3 1 3 3 3 3
1 3
18 3 3 1 3 3 0 3 1 0 2 0 0 1 3 3 1 3 3
14 3 0 3 0 1 3 3 0 1 3 3 1 3 0
19 3 0 1 2 1 3 2 0 2 1 1 0 1 0 1 0 1 0 0
3 3 3 0
5 3 3 1 0 1
7 3 3 2 3 0 1 3
9 3 3 1 3 3 0 1 3 3
3 3 0 3
6 3 0 3 0 3 0
7 3 1 3 0 0 1 3
2 3 3
17 3 0 3 1 3 0 3 0 1 2 1 0 2 2 0 3 0
6 3 1 1 3 1 3
4 3 0 2 3
4 3 0 3 0
1 3
4 3 0 2 3
4 3 1 3 0
2 3 3
13 3 0 3 1 2 1 1 3 3 3 3 0 3
1 3
2 3 0
6 3 0 3 0 0 3
13 3 0 3 1 0 1 2 3 3 1 3 3 3
4 3 1 3 0
18 3 0 3 1 3 3 1 3 2 3 1 1 1 1 1 1 1 1
6 3 1 3 1 3 0
5 3 1 3 3 0
6 3 1 3 0 1 0
12 3 3 1 3 3 0 3 1 3 2 0 3
3 3 0 3
3 3 1 2
15 3 1 1 3 3 0 0 3 0 1 2 3 0 0 0
9 3 0 3 1 3 0 3 1 3
2 3 3
2 3 3
8 3 1 1 3 0 0 1 3
4 3 0 2 3
12 3 0 2 3 0 1 2 1 3 0 2 1
6 3 3 1 3 3 3
8 3 0 3 0 2 0 3 0
7 3 0 3 0 0 1 2
6 3 1 3 1 3 3
5 3 0 0 2 3
3 3 0 3
7 3 0 3 1 2 2 3
12 3 0 3 0 3 0 3 3 1 3 3 3
19 3 0 1 3 3 1 0 1 2 1 2 0 3 0 3 0 1 0 3
9 3 0 3 1 3 2 0 3 0
3 3 1 3
15 3 0 3 0 3 1 3 3 0 2 3 2 3 0 3
7 3 0 3 0 1 3 3
5 3 0 2 1 3
2 3 1
6 3 3 1 3 3 3
8 3 3 0 0 3 3 0 3
2 3 3
5 3 1 3 0 1
15 3 3 1 1 1 1 1 1 1 1 1 1 3 1 3
22 3 0 2 3 0 0 0 1 1 2 1 2 3 1 0 1 3 3 0 2 0 3
4 3 3 3 2
3 3 3 3
3 3 1 3
3 3 3 2
11 3 0 3 1 2 2 3 1 3 3 2
4 3 3 3 0
4 3 3 3 2
36 3 0 1 3 3 0 2 3 3 1 3 0 2 0 2 3 0 1 3 3 3 3 0 1 1 0 0 1 3 3 3 1 1 0 1 3
2 3 1
11 3 0 3 0 1 2 3 0 3 0 1
8 3 1 3 0 1 1 2 0
3 3 0 3
7 3 0 3 1 2 0 3
4 3 1 3 1
7 3 0 3 1 0 1 0
2 3 3
5 3 0 3 1 2
3 3 1 3
6 3 0 2 3 1 3
1 3
18 3 1 1 0 3 3 3 3 0 2 1 0 2 3 1 2 3 1
5 3 0 2 1 3
14 3 3 1 3 3 3 0 3 3 0 1 0 3 1
6 3 1 1 3 0 1
11 3 3 1 3 3 3 0 2 2 0 3
1 3
3 3 1 2
21 3 3 2 0 2 0 2 3 1 3 3 0 3 1 2 3 0 1 2 1 3
4 3 3 0 2
3 3 0 3
12 3 1 3 0 2 3 2 1 1 2 1 3
10 3 1 3 1 3 3 3 1 0 3
19 3 0 3 1 2 3 0 0 0 2 0 3 0 1 3 3 0 1 2
13 3 3 0 1 2 3 1 3 3 1 3 0 2
2 3 3
8 3 3 2 1 3 3 1 3
3 3 0 3
16 3 0 1 1 3 3 3 3 3 3 3 0 1 3 3 3
1 3
2 3 3
3 3 1 2
1 3
8 3 0 3 0 1 3 3 3
17 3 3 3 2 3 0 2 2 2 3 0 2 0 3 0 1 3
6 3 0 1 0 0 3
7 3 3 1 3 3 0 3
3 3 3 0
3 3 3 1
3 3 1 3
14 3 0 3 3 0 1 2 3 1 3 1 0 3 0
7 3 0 3 1 2 3 0
7 3 0 3 1 3 0 2
24 3 0 3 1 2 2 0 2 3 3 1 1 3 3 0 3 1 3 3 0 1 3 1 2
47 3 0 2 3 1 3 2 1 2 0 3 1 3 1 3 1 1 1 1 1 1 3 0 1 3 3 3 1 1 1 1 3 1 3 0 0 2 0 3 1 3 0 1 3 3 0 1
6 3 3 1 2 3 0
3 3 0 3
4 3 3 0 2
21 3 3 0 2 1 1 3 3 1 1 3 1 3 3 0 3 1 3 3 2 1
3 3 0 3
3 3 3 0
3 3 1 3
9 3 0 3 1 2 1 0 3 1
9 3 0 3 0 1 3 3 1 3
4 3 1 3 0
9 3 1 1 1 3 3 3 0 2
11 3 0 3 1 0 1 2 3 3 0 0
6 3 0 3 0 2 0
3 3 0 3
3 3 3 0
3 3 0 3
15 3 3 1 0 1 3 3 1 1 1 3 1 3 0 2
8 3 3 0 0 0 3 3 3
4 3 0 3 3
5 3 0 3 3 0
3 3 3 0
3 3 1 3
7 3 0 3 1 2 1 3
7 3 0 3 2 0 3 0
1 3
9 3 3 3 0 3 3 3 3 0
6 3 3 0 0 1 3
6 3 0 3 0 0 1
1 3
12 3 0 3 0 3 0 1 3 3 1 3 2
2 3 3
2 3 3
5 3 3 1 1 0
6 3 3 1 2 1 1
2 3 3
6 3 0 3 1 3 0
25 3 3 0 2 0 1 0 2 3 1 2 2 0 3 0 3 0 3 1 2 1 1 1 3 1
6 3 3 0 3 0 3
1 3
12 3 3 0 1 1 0 2 0 2 3 0 0
8 3 3 0 3 1 2 0 2
10 3 0 3 0 2 0 1 3 1 0
6 3 0 3 2 0 3
4 3 0 3 0
4 3 1 1 3
6 3 0 3 1 2 3
6 3 3 3 1 1 3
9 3 1 2 0 1 2 3 0 1
7 3 3 1 3 3 1 3
5 3 3 0 0 0
8 3 1 2 3 0 2 1 2
3 3 0 3
3 3 3 1
3 3 1 3
10 3 0 3 0 2 0 0 2 0 3
4 3 3 0 0
9 3 3 1 3 3 2 0 3 0
1 3
4 3 3 1 3
3 3 1 3
4 3 3 0 0
3 3 0 3
2 3 3
5 3 3 0 1 0
6 3 1 1 1 3 3
8 3 0 3 0 1 0 1 3
6 3 3 1 3 3 1
5 3 2 0 1 3
7 3 0 3 1 3 1 3
1 3
2 3 3
23 3 0 3 3 3 3 2 1 0 2 0 3 0 2 0 3 0 1 3 3 0 2 0
5 3 3 3 3 3
3 3 3 0
9 3 0 3 0 1 0 0 2 3
6 3 3 0 0 3 0
6 3 0 2 3 3 0
28 3 1 2 1 3 0 0 1 0 0 1 3 3 3 0 0 3 1 3 1 1 3 2 0 1 1 1 0
8 3 0 3 1 3 1 2 3
4 3 0 3 3
9 3 3 0 0 3 3 0 0 2
7 3 0 3 0 2 0 3
3 3 3 1
3 3 0 3
3 3 1 3
4 3 0 2 3
5 3 3 1 0 2
6 3 0 3 1 3 0
3 3 3 0
5 3 0 3 3 3
1 3
1 3
10 3 3 2 0 2 3 1 2 0 3
21 3 0 3 1 3 0 3 1 2 1 1 2 3 1 1 1 2 0 2 1 3
3 3 3 0
13 3 0 3 0 3 0 1 3 3 3 1 3 0
2 3 3
10 3 0 1 3 3 1 3 0 1 0
2 3 3
3 3 0 3
5 3 1 1 3 1
9 3 0 3 1 2 3 1 3 3
23 3 0 3 0 1 2 1 2 0 3 3 1 3 3 0 3 0 3 0 3 1 2 3
3 3 0 2
1 3
6 3 3 0 2 1 0
4 3 2 0 3
7 3 3 2 1 3 3 0
6 3 1 1 3 0 1
4 3 1 3 0
5 3 0 0 0 3
3 3 1 3
2 3 1
3 3 3 0
7 3 0 3 1 3 0 1
4 3 0 3 0
2 3 3
3 3 0 3
5 3 2 0 3 0
2 3 3
6 3 0 1 2 3 3
3 3 1 2
6 3 0 3 0 2 3
8 3 3 1 3 3 1 0 2
12 3 0 2 3 0 0 0 2 3 2 1 0
9 3 0 3 0 1 3 3 1 3
6 3 0 2 1 1 3
7 3 0 2 2 0 3 0
8 3 0 3 1 0 2 1 3
2 3 3
8 3 1 1 3 0 2 3 0
5 3 3 1 3 3
3 3 3 2
2 3 0
12 3 0 3 0 1 3 3 0 3 0 3 0
2 3 0
3 3 3 2
2 3 1
4 3 0 3 0
13 3 3 0 0 1 3 0 1 3 2 0 3 0
14 3 0 2 0 1 3 1 1 1 1 2 1 3 0
9 3 0 3 2 3 3 1 1 3
2 3 0
3 3 0 3
3 3 3 0
21 3 3 2 1 0 1 3 3 1 2 1 1 1 2 0 3 0 3 3 0 2
5 3 0 3 1 2
4 3 3 0 2
21 3 3 1 3 3 0 3 0 1 3 3 3 0 0 2 2 3 0 1 2 3
7 3 1 1 1 1 1 3
4 3 1 3 0
18 3 0 3 3 1 0 0 3 1 1 0 1 0 0 2 1 1 0
5 3 3 0 1 1
15 3 1 3 0 0 1 3 0 2 0 3 1 2 3 0
4 3 0 2 3
8 3 3 0 2 0 2 1 3
3 3 0 3
11 3 3 1 1 2 0 2 3 1 2 1
17 3 0 2 3 1 3 3 0 3 0 1 1 1 2 1 3 0
2 3 3
18 3 3 1 3 3 0 1 1 2 3 1 3 3 0 0 1 1 3
5 3 3 1 3 3
13 3 3 0 1 1 2 0 3 0 3 0 0 3
16 3 1 2 1 3 3 3 3 0 0 1 1 3 1 3 0
13 3 3 3 3 0 1 0 1 2 0 1 3 0
8 3 3 1 3 3 1 3 0
4 3 3 0 2
12 3 0 3 1 3 1 3 0 2 2 0 3
15 3 0 3 0 1 1 3 3 0 2 1 0 0 3 2
5 3 0 1 1 1
5 3 3 2 1 0
5 3 1 3 0 2
13 3 0 3 0 1 3 3 3 2 0 2 0 3
26 3 3 0 3 3 3 0 1 1 1 1 1 0 2 0 3 0 2 0 0 2 1 1 3 3 3
2 3 3
9 3 2 0 3 1 3 3 0 3
2 3 3
9 3 0 3 1 3 3 2 0 0
3 3 3 0
16 3 0 1 3 3 3 0 2 0 3 0 2 1 1 0 2
14 3 0 3 0 1 3 3 0 3 0 2 3 0 2
9 3 3 2 3 1 0 3 2 2
5 3 3 0 0 0
3 3 0 3
2 3 1
3 3 1 3
2 3 3
6 3 3 1 3 3 1
4 3 0 3 0
2 3 0
2 3 3
9 3 1 3 0 2 0 3 1 3
16 3 0 3 3 3 1 2 2 0 3 1 3 0 3 3 3
9 3 0 3 0 1 3 3 0 1
3 3 3 0
2 3 3
9 3 3 0 0 1 1 3 0 0
2 3 3
3 3 0 3
3 3 3 1
4 3 2 0 3
4 3 3 0 0
5 3 0 3 0 2
2 3 3
8 3 1 1 1 1 1 1 1
7 3 0 3 0 2 0 3
16 3 0 3 0 3 0 1 0 0 1 3 3 3 0 2 3
7 3 1 3 0 1 2 3
2 3 3
9 3 0 3 1 2 3 0 0 0
11 3 0 3 0 3 1 3 1 3 0 2
2 3 3
2 3 2
12 3 0 3 1 2 1 2 0 3 3 0 0
2 3 3
7 3 3 0 2 3 2 0
4 3 3 2 0
10 3 3 1 3 3 0 1 0 3 3
13 3 0 3 0 1 2 0 2 1 3 3 2 3
1 3
3 3 1 2
1 3
2 3 2
5 3 3 1 3 3
3 3 1 3
28 3 1 1 3 1 2 0 2 0 1 3 3 0 1 2 3 0 0 1 3 1 1 1 3 3 2 2 3
8 3 0 3 0 0 3 0 2
19 3 3 0 2 3 1 3 3 1 0 1 2 3 0 0 3 3 0 3
17 3 0 3 3 0 1 3 2 1 2 0 3 0 3 1 2 3
9 3 1 3 1 1 3 3 3 1
6 3 0 3 0 1 3
30 3 1 2 3 0 3 3 0 3 0 3 3 1 3 3 0 2 0 3 1 3 3 1 0 1 0 0 0 2 0
1 3
1 3
5 3 1 0 1 3
5 3 3 0 0 0
3 3 1 3
12 3 1 2 1 3 3 3 1 3 3 1 3
5 3 3 1 0 3
6 3 3 2 0 0 0
3 3 1 3
10 3 3 1 1 1 1 1 0 1 1
3 3 3 2
2 3 3
3 3 3 0
21 3 3 1 3 2 0 0 1 1 1 1 1 2 0 3 1 2 3 1 2 3
15 3 1 3 0 2 0 3 1 0 1 3 3 0 1 0
11 3 0 2 0 0 1 2 3 1 3 0
9 3 3 0 1 1 3 2 0 3
9 3 3 1 3 3 1 3 0 3
8 3 3 3 1 3 3 1 3
3 3 0 3
7 3 3 1 1 1 2 0
16 3 1 1 3 0 1 3 2 1 2 0 3 0 1 2 3
2 3 3
1 3
7 3 0 3 1 3 0 2
17 3 3 1 3 3 3 0 1 1 0 2 0 3 1 2 0 3
18 3 0 1 2 2 3 1 3 3 0 3 2 0 3 1 3 3 0
12 3 0 3 1 2 1 1 3 2 1 1 3
3 3 0 3
1 3
8 3 3 2 0 1 1 1 0
5 3 0 3 3 0
3 3 0 3
2 3 3
6 3 3 1 3 3 3
4 3 1 1 3
7 3 0 1 3 3 3 0
3 3 1 3
5 3 1 0 3 3
7 3 0 0 3 2 1 3
9 3 3 0 2 1 1 3 3 3
2 3 3
7 3 0 3 1 2 1 0
2 3 3
18 3 3 2 0 2 3 1 2 1 2 3 1 3 3 0 3 3 1
12 3 3 1 3 3 0 1 3 3 3 0 2
1 3
4 3 1 3 0
10 3 3 0 2 1 1 3 0 3 3
2 3 3
2 3 3
11 3 0 3 0 3 3 1 2 0 2 1
8 3 0 3 0 1 2 1 0
12 3 1 3 0 1 1 1 1 2 3 1 0
3 3 1 3
17 3 0 0 2 3 1 3 2 0 0 2 1 2 0 2 0 3
17 3 3 1 3 3 3 3 3 3 1 0 1 3 3 0 1 2
11 3 0 3 2 0 1 3 1 0 3 0
11 3 3 1 1 1 2 1 3 0 1 0
2 3 3
1 3
3 3 3 1
11 3 3 1 3 3 0 3 0 1 2 3
7 3 0 3 1 3 1 3
5 3 3 0 1 0
16 3 0 3 1 2 1 1 3 2 2 0 3 0 2 0 3
9 3 0 3 1 3 0 3 1 3
18 3 0 3 0 1 3 3 1 2 3 1 2 1 1 1 1 0 1
7 3 0 3 1 3 3 0
2 3 3
7 3 0 3 0 1 2 3
4 3 3 0 0
6 3 0 3 0 1 0
2 3 3
2 3 3
3 3 1 3
7 3 0 3 1 2 1 1
6 3 1 3 0 0 3
5 3 0 3 0 3
4 3 0 3 0
3 3 3 3
1 3
13 3 2 0 3 0 2 0 3 0 3 0 2 3
5 3 1 3 1 0
14 3 0 3 0 2 3 2 3 0 0 2 0 0 2
12 3 0 3 0 3 0 1 3 3 0 2 3
9 3 1 2 0 0 3 0 0 2
17 3 0 3 1 2 2 0 3 0 1 1 3 3 1 3 0 3
5 3 2 0 3 0
26 3 3 0 0 0 1 3 3 3 1 3 0 3 0 1 3 3 1 2 1 2 1 0 1 1 3
1 3
7 3 3 3 0 2 0 3
4 3 0 2 3
3 3 1 3
6 3 3 0 0 1 3
3 3 0 3
1 3
9 3 3 1 3 3 3 1 0 2
4 3 3 0 2
1 3
15 3 1 3 2 0 0 1 3 0 0 3 3 0 3 0
5 3 0 3 3 2
10 3 0 3 3 1 3 3 3 2 0
8 3 0 3 1 2 1 3 1
7 3 0 3 1 3 0 3
35 3 0 3 0 0 1 2 2 0 2 3 0 0 0 3 3 3 0 1 1 1 3 3 3 0 1 3 3 3 0 0 0 1 3 3
5 3 0 1 0 3
3 3 3 0
13 3 0 3 3 0 0 3 3 3 3 3 1 3
13 3 0 3 1 3 3 0 1 2 3 2 0 2
2 3 3
8 3 1 1 3 0 0 0 1
5 3 0 3 3 0
7 3 0 2 3 1 3 3
17 3 1 0 3 3 0 0 3 0 2 1 1 1 1 3 1 3
1 3
5 3 3 0 2 3
2 3 1
7 3 3 3 0 1 0 1
4 3 3 1 0
6 3 3 0 2 0 3
7 3 0 1 1 3 3 3
12 3 3 0 1 2 3 0 2 3 1 3 3
23 3 1 0 3 3 0 1 3 3 0 3 0 1 3 3 1 2 3 0 1 2 0 3
3 3 0 3
10 3 1 3 0 1 1 2 0 3 3
4 3 0 3 0
9 3 1 3 2 1 0 2 3 2
19 3 0 2 3 1 3 3 1 2 1 3 0 2 1 1 1 1 1 1
4 3 0 1 0
21 3 1 3 1 1 3 2 1 2 0 3 1 0 1 3 3 1 2 0 3 0
32 3 0 3 1 0 1 0 1 2 3 0 2 0 3 0 2 3 0 2 0 3 0 1 2 2 0 3 0 1 3 3 0
4 3 3 0 0
5 3 2 0 3 0
5 3 3 1 3 3
5 3 3 3 2 0
7 3 1 1 1 3 3 2
6 3 3 1 3 3 3
2 3 3
8 3 3 1 3 3 0 0 1
27 3 0 3 0 1 3 3 0 1 3 3 1 3 3 1 3 3 0 1 0 1 3 0 2 2 0 3
10 3 0 3 0 1 3 3 0 3 0
3 3 3 0
2 3 3
9 3 1 3 1 3 3 1 3 3
5 3 1 3 0 0
2 3 3
3 3 3 2
6 3 3 2 0 3 3
2 3 2
2 3 3
7 3 3 1 1 1 1 2
24 3 1 3 0 1 3 1 3 3 3 0 3 0 3 0 1 2 2 0 3 0 1 0 3
2 3 3
21 3 0 3 0 3 2 0 1 3 0 0 3 3 2 0 1 1 1 2 0 1
8 3 3 1 3 3 1 3 2
2 3 3
4 3 2 0 3
4 3 0 2 3
3 3 0 3
3 3 3 3
8 3 1 1 3 0 2 1 3
11 3 3 0 1 1 1 0 2 1 1 2
4 3 0 2 3
1 3
4 3 0 3 3
1 3
3 3 0 3
3 3 0 3
12 3 0 3 1 0 1 2 3 3 0 0 0
11 3 0 3 0 3 3 1 3 3 0 2
7 3 3 1 2 3 0 1
3 3 1 3
6 3 0 3 1 3 3
6 3 1 1 3 0 0
28 3 0 1 0 3 3 0 1 3 1 3 3 1 3 0 2 0 2 3 0 1 1 1 3 1 1 2 3
3 3 1 3
4 3 0 3 0
8 3 0 3 1 1 3 1 3
4 3 0 1 2
1 3
3 3 1 3
5 3 3 2 0 0
9 3 1 1 3 0 2 3 1 0
18 3 0 3 0 3 0 1 2 1 0 3 3 0 3 3 0 1 0
13 3 1 3 0 1 1 1 0 0 0 1 3 3
3 3 0 3
7 3 0 1 3 3 1 3
11 3 3 0 1 0 0 1 2 1 1 3
15 3 0 3 0 3 1 0 1 0 0 2 2 2 3 0
26 3 0 3 0 1 3 3 0 0 1 1 2 3 1 2 1 0 1 1 3 0 2 0 3 1 2
3 3 0 2
7 3 0 3 1 3 1 3
6 3 0 3 3 0 0
2 3 3
3 3 3 0
3 3 0 3
1 3
4 3 0 0 0
3 3 0 3
5 3 3 1 1 3
9 3 0 3 0 2 2 2 3 0
7 3 2 0 3 0 1 3
6 3 3 2 0 0 0
2 3 3
3 3 3 0
3 3 0 2
8 3 0 3 0 1 2 0 0
23 3 0 3 0 3 0 1 1 3 3 2 3 1 1 3 1 3 0 2 3 1 3 3
3 3 0 3
9 3 0 3 0 1 2 0 3 0
3 3 3 0
19 3 0 2 1 0 1 1 0 1 3 3 0 3 1 0 2 2 1 3
15 3 0 3 0 1 2 1 3 0 0 3 0 0 0 0
3 3 1 2
1 3
8 3 1 0 3 3 1 3 2
6 3 1 3 1 3 3
9 3 1 1 3 1 3 1 3 3
14 3 0 3 0 1 2 0 0 3 1 3 3 0 3
9 3 1 0 0 0 2 1 3 2
14 3 3 1 0 0 1 3 0 2 0 2 1 3 1
7 3 3 1 3 3 3 3
3 3 0 3
5 3 3 1 3 1
5 3 3 1 0 0
5 3 3 0 0 0
3 3 3 0
1 3
4 3 1 3 0
5 3 1 3 0 2
4 3 3 2 0
6 3 0 3 0 1 2
4 3 1 1 3
7 3 0 3 1 0 2 1
4 3 1 3 0
5 3 3 1 3 3
9 3 3 1 0 3 1 1 0 0
9 3 0 3 0 1 2 2 0 1
2 3 3
6 3 0 3 1 3 3
15 3 1 3 0 1 1 0 1 2 2 0 3 0 1 0
3 3 1 3
20 3 0 2 2 3 0 2 3 2 1 3 1 3 3 3 3 3 1 0 3
6 3 3 3 2 1 3
8 3 1 3 0 2 1 1 2
17 3 3 0 1 3 3 3 3 0 3 1 0 1 3 3 3 2
3 3 0 3
15 3 3 0 1 2 3 1 3 3 1 3 0 0 1 3
1 3
3 3 1 1
1 3
5 3 3 0 0 3
3 3 0 3
1 3
2 3 3
4 3 0 2 3
11 3 3 0 1 1 3 3 3 3 0 2
11 3 3 1 3 0 2 2 2 3 0 0
1 3
19 3 3 2 0 2 1 3 1 3 3 3 1 3 3 0 2 2 2 3
17 3 0 3 3 3 0 2 0 3 0 0 2 3 2 0 1 3
5 3 0 3 1 0
7 3 3 1 2 3 1 3
3 3 1 2
12 3 0 3 1 0 1 1 3 2 1 1 3
13 3 3 0 2 1 2 0 0 1 3 0 0 3
30 3 3 1 3 3 0 3 0 1 3 3 3 0 2 0 3 0 1 0 1 2 3 0 3 0 1 3 3 0 2
2 3 3
9 3 3 1 3 1 1 1 2 0
2 3 3
4 3 1 3 0
23 3 0 1 3 3 0 3 0 1 3 3 3 0 1 2 3 0 1 1 1 2 0 3
7 3 2 0 3 0 0 3
13 3 3 0 1 2 3 1 3 3 0 3 3 1
8 3 1 1 3 3 1 3 2
10 3 3 3 1 3 3 0 1 3 3
3 3 1 3
8 3 0 3 3 0 3 3 1
4 3 3 0 1
1 3
3 3 3 0
1 3
3 3 0 3
3 3 3 3
2 3 3
5 3 3 0 1 0
2 3 3
29 3 0 2 3 3 3 3 3 3 3 0 1 0 1 3 3 3 1 3 3 3 1 2 1 1 1 2 1 3
4 3 1 2 3
3 3 1 2
5 3 1 3 0 0
7 3 2 0 3 0 1 1
5 3 0 2 2 3
16 3 3 0 2 0 3 0 1 3 3 3 1 3 2 1 1
2 3 3
8 3 3 0 1 2 1 3 0
14 3 0 3 3 1 3 3 0 2 3 0 2 0 2
5 3 3 1 0 0
2 3 3
3 3 0 3
6 3 0 1 0 1 3
6 3 0 2 1 3 0
3 3 3 2
2 3 3
5 3 3 0 0 0
10 3 0 3 0 3 1 3 0 2 3
11 3 3 3 3 2 1 1 2 0 3 0
12 3 3 1 3 3 0 1 1 3 3 0 3
6 3 0 3 1 2 3
9 3 3 0 0 3 3 0 3 1
2 3 3
3 3 1 3
8 3 0 3 0 1 2 3 3
9 3 0 3 0 3 0 0 2 2
7 3 0 3 1 2 0 3
10 3 3 1 3 3 0 3 1 3 3
3 3 3 0
33 3 0 1 3 3 1 3 0 3 0 3 0 3 1 3 1 3 3 2 0 3 0 1 1 1 3 1 2 1 3 0 1 0
4 3 0 2 3
12 3 0 3 3 3 0 3 0 1 3 3 3
8 3 0 3 1 2 1 1 3
2 3 3
29 3 0 3 3 0 1 3 3 3 3 3 0 1 3 3 3 3 1 0 1 3 1 2 1 1 3 3 3 0
3 3 1 3
3 3 1 3
8 3 1 2 0 1 2 3 0
1 3
2 3 3
21 3 1 3 0 1 0 1 3 3 3 1 2 1 3 2 1 1 1 3 1 3
4 3 1 1 3
15 3 0 3 0 1 2 2 0 0 0 0 3 3 3 3
4 3 1 1 3
10 3 0 3 0 1 0 1 3 3 0
4 3 0 2 3
4 3 0 3 3
4 3 0 3 3
1 3
4 3 1 3 2
2 3 3
2 3 3
3 3 0 3
2 3 3
2 3 3
2 3 3
6 3 1 3 3 1 3
2 3 3
8 3 0 3 1 2 3 0 0
13 3 0 0 1 1 3 1 3 3 3 1 1 1
3 3 1 3
6 3 0 0 3 0 2
2 3 3
4 3 0 3 3
26 3 1 2 1 1 3 3 0 3 0 3 0 3 0 3 0 3 0 2 3 0 0 1 3 0 2
2 3 0
2 3 3
17 3 3 3 1 1 3 2 1 1 3 0 1 3 3 1 3 3
3 3 0 3
1 3
6 3 0 3 0 2 1
7 3 0 3 0 3 0 3
2 3 1
5 3 0 3 0 1
11 3 1 3 0 0 1 1 3 1 2 1
3 3 1 3
2 3 0
2 3 3
2 3 0
8 3 0 3 0 1 3 3 3
1 3
4 3 3 3 0
10 3 3 0 1 1 1 1 2 1 3
8 3 0 3 2 3 1 3 3
3 3 1 3
9 3 3 1 2 2 3 1 3 3
4 3 2 0 3
12 3 0 3 0 1 3 3 3 0 0 3 0
12 3 3 0 1 1 2 3 1 3 3 0 3
11 3 0 3 0 1 3 3 0 1 3 3
8 3 1 3 1 3 1 3 0
13 3 3 2 0 0 3 3 3 3 3 2 0 3
3 3 0 3
4 3 0 3 3
1 3
11 3 0 3 1 1 1 1 1 1 1 1
7 3 0 3 0 1 3 3
25 3 0 3 0 1 3 1 2 1 3 0 1 1 2 1 0 1 3 3 3 2 0 3 0 2
26 3 3 1 3 3 1 1 1 3 1 3 3 3 1 3 3 3 1 3 3 1 3 0 2 0 3
3 3 1 2
6 3 0 3 1 3 0
5 3 1 3 1 3
10 3 1 0 1 1 3 0 2 1 2
8 3 0 3 1 2 0 1 3
3 3 3 0
8 3 0 3 3 0 0 3 3
3 3 3 0
6 3 3 0 3 3 3
5 3 0 3 1 3
1 3
12 3 0 3 1 2 3 0 2 0 3 0 3
6 3 1 0 3 1 3
4 3 0 2 3
3 3 0 3
5 3 0 3 0 2
1 3
12 3 3 2 1 2 3 0 3 0 3 3 3
2 3 3
2 3 3
16 3 0 3 0 1 0 2 0 0 2 3 1 3 2 0 0
10 3 1 3 0 1 3 1 0 3 0
5 3 3 1 3 3
1 3
12 3 0 3 0 1 3 3 0 2 3 1 2
9 3 0 3 0 0 1 2 0 3
4 3 0 2 3
2 3 3
1 3
2 3 3
2 3 3
6 3 0 3 0 3 0
4 3 0 3 3
19 3 3 0 2 0 1 0 1 2 2 0 3 3 3 1 1 0 0 1
1 3
2 3 3
3 3 0 3
14 3 0 3 1 3 0 3 0 1 3 3 0 2 1
4 3 3 0 0
8 3 0 3 0 3 3 0 0
16 3 0 2 3 0 2 0 3 1 1 1 1 1 1 0 1
2 3 3
17 3 1 1 1 1 1 1 1 1 1 1 1 2 3 0 0 1
3 3 3 0
4 3 0 2 3
9 3 0 3 1 2 2 0 2 3
13 3 0 3 0 1 0 1 0 1 3 3 1 3
5 3 0 1 3 3
13 3 0 3 1 1 3 0 1 1 2 3 3 2
3 3 3 2
11 3 3 0 1 1 2 0 1 2 3 1
12 3 0 3 1 2 0 0 3 0 0 1 3
12 3 3 0 1 1 2 3 1 3 0 2 3
5 3 3 1 3 3
16 3 3 0 2 1 3 2 0 2 0 1 2 1 0 3 2
6 3 3 2 3 2 2
14 3 1 3 3 3 0 3 0 2 3 0 0 0 2
1 3
4 3 1 3 0
16 3 3 1 1 1 1 1 1 3 1 3 1 3 3 0 2
3 3 3 3
6 3 3 0 0 0 1
3 3 0 3
6 3 0 3 0 2 2
3 3 0 3
5 3 0 3 3 3
14 3 1 3 0 2 1 0 3 3 0 2 1 1 3
3 3 0 3
6 3 3 1 3 3 1
6 3 2 1 0 0 1
1 3
2 3 0
3 3 0 1
1 3
13 3 3 3 1 3 3 3 3 1 3 3 0 2
3 3 0 1
3 3 1 2
6 3 0 3 0 3 0
1 3
4 3 0 2 3
3 3 1 3
3 3 1 3
2 3 3
5 3 1 1 3 0
8 3 0 3 0 1 2 0 2
8 3 1 2 1 1 3 0 3
5 3 3 0 0 0
2 3 3
10 3 3 1 2 3 3 0 1 1 0
7 3 3 0 2 0 0 0
3 3 1 3
10 3 0 3 1 2 1 1 1 1 0
2 3 3
14 3 0 3 0 1 0 1 3 3 0 1 0 0 2
11 3 0 1 2 1 2 0 3 1 2 3
7 3 0 3 1 2 0 3
2 3 3
11 3 0 3 0 3 1 3 1 1 3 0
11 3 0 3 0 2 3 0 3 0 1 0
5 3 0 3 1 0
1 3
2 3 3
11 3 3 1 3 3 0 3 0 1 3 2
2 3 3
26 3 3 0 2 1 1 2 3 0 0 1 3 0 2 3 3 0 1 2 1 1 3 3 2 0 0
22 3 1 3 1 3 2 1 3 1 3 2 1 1 1 1 1 1 2 0 3 0 2
3 3 1 3
11 3 3 0 1 3 0 1 0 3 1 0
3 3 1 3
3 3 0 3
11 3 3 1 3 3 0 3 1 2 1 0
3 3 1 3
3 3 0 3
5 3 3 0 3 3
4 3 3 2 0
3 3 1 3
5 3 1 3 0 0
7 3 3 1 3 3 0 2
5 3 2 0 1 3
8 3 1 3 0 1 3 1 1
18 3 0 3 0 1 3 3 0 3 1 0 1 3 3 0 2 3 3
4 3 1 3 0
6 3 2 0 1 3 0
13 3 0 3 0 3 0 1 3 2 0 1 3 3
2 3 3
1 3
2 3 3
2 3 2
4 3 1 3 0
8 3 3 2 3 0 2 0 3
5 3 1 1 3 3
15 3 0 3 0 0 0 1 2 0 3 3 1 1 1 3
3 3 1 3
3 3 3 2
7 3 3 0 2 1 3 0
4 3 1 0 3
5 3 3 0 1 1
5 3 0 0 3 2
9 3 0 1 1 1 3 2 3 0
3 3 0 1
1 3
9 3 0 3 0 1 0 1 2 3
6 3 0 3 3 0 2
2 3 3
14 3 0 2 3 1 0 1 1 1 1 1 1 0 1
6 3 0 3 1 3 3
2 3 0
54 3 3 0 2 1 1 1 1 3 3 2 1 3 2 2 0 3 3 0 2 0 3 1 0 1 3 3 3 1 1 1 1 1 1 1 2 0 3 1 2 1 3 3 1 1 3 0 2 0 3 1 3 3 0
2 3 1
15 3 0 0 2 2 1 3 0 0 1 3 0 2 0 2
5 3 3 3 2 0
2 3 3
5 3 0 3 0 3
9 3 1 3 1 3 0 1 2 0
3 3 0 2
7 3 3 1 2 3 3 0
14 3 1 3 1 3 3 1 2 1 0 1 1 0 3
5 3 0 3 1 0
4 3 3 0 2
3 3 1 2
5 3 3 0 0 3
8 3 0 2 1 1 3 3 2
2 3 3
8 3 0 3 0 1 3 3 0
4 3 3 0 0
2 3 3
8 3 3 1 3 3 0 2 3
6 3 1 3 0 0 0
3 3 0 3
3 3 0 3
3 3 1 3
2 3 3
14 3 1 1 3 1 3 3 3 0 2 1 1 0 0
8 3 3 0 1 1 1 2 0
17 3 0 2 3 1 3 3 0 3 0 3 3 0 1 1 1 0
6 3 0 3 3 3 1
12 3 0 3 1 3 0 3 1 3 1 2 0
3 3 3 0
4 3 1 3 3
2 3 3
3 3 1 3
8 3 0 3 0 1 3 3 0
11 3 0 3 0 1 2 1 3 2 1 0
8 3 1 3 0 1 1 0 1
3 3 0 3
4 3 3 0 0
2 3 3
6 3 3 0 2 0 3
10 3 1 3 1 1 3 2 3 0 2
2 3 3
16 3 3 0 2 1 1 3 3 0 2 0 1 3 1 3 2
5 3 3 0 1 0
3 3 0 1
3 3 1 3
6 3 0 3 0 3 3
13 3 0 3 0 1 2 0 1 1 1 3 0 2
12 3 3 0 2 3 1 3 0 3 1 2 1
6 3 3 0 3 3 0
7 3 3 0 1 0 1 1
1 3
2 3 3
9 3 1 0 3 1 2 2 0 3
2 3 3
7 3 3 0 2 1 3 2
1 3
11 3 3 0 0 3 3 3 3 3 1 3
3 3 0 3
6 3 0 3 0 1 0
5 3 3 0 1 0
5 3 3 1 3 0
2 3 3
8 3 0 3 1 3 0 1 0
3 3 0 3
13 3 0 2 1 1 2 1 2 3 1 2 1 3
3 3 1 3
10 3 1 1 3 0 1 2 3 1 0
2 3 3
3 3 3 0
3 3 0 3
2 3 3
14 3 0 3 0 1 3 3 3 3 1 3 3 3 0
8 3 0 3 0 1 0 1 3
36 3 0 3 2 0 3 0 1 1 2 3 1 3 3 3 0 0 1 1 3 0 2 0 3 0 3 1 3 0 3 0 3 0 1 0 0
3 3 3 0
6 3 0 3 0 1 2
3 3 1 3
3 3 3 2
4 3 1 3 0
10 3 0 3 1 3 0 3 0 1 2
10 3 3 0 0 0 3 1 3 2 1
27 3 3 0 0 3 3 1 1 1 1 0 1 0 2 0 1 2 0 3 1 3 3 3 1 0 0 1
2 3 3
21 3 3 2 0 1 1 1 1 0 0 1 3 3 0 1 3 3 0 3 0 2
10 3 3 0 0 3 3 3 3 3 3
8 3 3 0 1 2 0 3 0
12 3 0 3 0 0 0 0 1 3 3 1 0
6 3 0 3 1 2 1
10 3 0 2 3 0 2 1 0 3 0
3 3 0 3
2 3 3
6 3 3 1 2 1 1
16 3 0 3 0 3 1 3 0 1 3 2 1 0 2 1 2
7 3 3 1 2 3 0 3
8 3 0 3 1 2 0 3 0
16 3 0 3 1 0 2 0 1 3 0 3 0 2 0 0 0
6 3 0 3 0 3 3
20 3 0 3 1 1 3 3 3 0 3 1 3 3 0 0 3 2 1 1 3
4 3 3 2 0
2 3 3
4 3 1 1 3
4 3 3 0 1
21 3 1 3 0 1 1 3 3 3 3 1 2 3 0 2 0 3 1 2 0 3
17 3 0 3 1 2 0 2 1 0 1 1 3 3 0 1 2 3
9 3 1 3 0 1 2 0 3 0
2 3 3
3 3 3 0
19 3 0 2 3 1 2 1 1 2 1 0 3 3 1 3 1 3 0 2
8 3 3 1 3 0 2 0 3
4 3 0 2 3
8 3 0 3 0 0 2 3 3
2 3 3
7 3 1 1 3 1 3 3
1 3
5 3 0 1 0 0
2 3 0
15 3 0 3 1 0 2 2 2 3 1 3 1 3 0 1
7 3 0 3 0 2 0 3
14 3 3 1 3 3 1 2 1 0 1 3 3 3 1
23 3 3 2 3 1 3 3 0 1 2 0 1 0 1 3 1 3 3 0 1 3 3 0
2 3 3
2 3 3
2 3 3
3 3 0 3
2 3 3
2 3 3
20 3 0 3 0 2 1 3 0 2 0 3 3 1 3 3 0 3 1 1 3
2 3 3
2 3 3
3 3 0 3
4 3 0 2 3
6 3 0 3 0 2 3
15 3 0 3 1 2 2 0 3 0 3 1 2 3 0 1
32 3 0 3 3 3 1 3 2 1 1 1 1 2 0 3 1 3 3 2 0 2 0 3 0 2 0 3 0 2 0 3 3
26 3 0 3 0 0 3 0 1 3 3 0 1 1 1 1 1 3 2 3 0 2 3 2 3 1 2
12 3 2 0 1 3 0 1 3 1 2 0 3
2 3 3
7 3 0 3 1 2 1 1
7 3 0 3 1 2 0 3
9 3 1 1 1 3 0 1 3 0
25 3 3 0 1 2 0 2 3 1 1 3 1 3 1 3 3 0 3 0 2 0 0 0 1 0
13 3 0 3 0 1 0 0 2 3 2 3 0 0
20 3 3 1 3 3 1 3 0 2 2 3 0 2 0 0 1 3 3 0 2
11 3 3 1 3 3 0 3 3 3 1 2
3 3 0 3
2 3 0
5 3 2 0 3 0
12 3 0 3 1 2 1 1 1 0 1 2 3
6 3 3 0 2 3 3
7 3 0 0 0 3 2 3
54 3 3 0 2 1 1 3 0 2 3 1 1 3 0 1 3 1 0 1 2 3 0 3 1 2 2 0 3 1 0 1 3 3 0 2 3 0 1 1 1 1 3 1 0 1 2 0 3 1 3 0 2 3 0
9 3 0 3 1 2 1 2 0 3
7 3 1 3 0 2 1 2
35 3 2 0 3 3 3 2 3 0 0 3 3 3 3 3 2 0 3 0 2 1 1 3 0 2 0 3 0 1 3 3 0 3 1 3
18 3 0 3 1 2 1 3 1 3 2 3 0 3 0 3 0 2 0
4 3 0 1 2
13 3 0 3 0 2 3 0 3 1 2 1 0 1
2 3 0
1 3
10 3 3 1 3 3 1 0 1 3 3
8 3 3 1 3 0 3 3 3
3 3 3 0
22 3 3 1 3 3 3 3 0 0 1 3 1 1 1 3 1 1 1 2 0 3 3
7 3 0 3 3 3 0 3
3 3 1 3
4 3 0 2 0
1 3
3 3 0 2
10 3 3 0 1 1 1 1 1 0 1
3 3 3 0
2 3 3
2 3 3
2 3 3
2 3 3
7 3 3 1 3 3 0 3
3 3 0 3
15 3 0 0 3 2 1 0 2 0 2 3 0 1 1 3
2 3 3
10 3 3 0 0 3 3 1 1 2 3
6 3 3 2 3 1 3
1 3
9 3 3 1 3 3 0 1 3 3
3 3 3 2
11 3 0 3 1 3 0 3 3 1 2 3
7 3 0 3 0 1 3 3
9 3 3 3 2 3 0 2 1 3
7 3 0 3 1 3 0 1
19 3 0 3 1 2 1 1 2 1 3 0 1 2 0 2 1 1 3 0
16 3 0 3 0 1 1 3 2 0 3 1 1 3 1 1 3
5 3 3 1 0 0
13 3 2 2 1 2 1 2 3 1 3 3 3 2
24 3 0 3 0 3 1 0 1 2 3 1 3 0 1 1 1 1 2 0 3 1 2 0 3
3 3 0 1
6 3 0 3 0 2 3
1 3
9 3 0 3 0 3 0 3 1 3
3 3 3 2
8 3 3 1 1 3 3 3 0
2 3 3
4 3 1 3 0
9 3 0 3 2 0 1 1 3 0
5 3 0 3 1 3
3 3 3 0
10 3 3 0 2 1 1 1 1 1 3
1 3
2 3 3
2 3 3
4 3 2 0 3
1 3
1 3
12 3 0 3 1 2 1 3 1 0 1 2 3
9 3 0 3 1 0 1 3 3 3
7 3 0 2 1 1 1 3
3 3 0 3
2 3 3
10 3 3 3 2 0 2 0 3 1 0
17 3 0 3 0 3 3 1 3 3 0 2 3 3 1 3 0 1
20 3 0 3 0 1 1 3 0 3 3 1 1 3 1 3 2 1 1 1 3
3 3 0 3
24 3 3 0 2 1 1 1 3 0 0 1 2 3 0 1 3 2 0 0 2 3 0 1 1
11 3 3 2 0 3 3 3 0 0 0 3
5 3 1 3 0 2
4 3 3 0 2
12 3 2 0 3 0 1 1 1 1 2 0 3
1 3
3 3 1 1
11 3 1 3 0 2 0 3 1 0 2 3
2 3 3
2 3 0
3 3 0 1
2 3 3
2 3 3
11 3 0 3 0 1 3 3 1 3 3 0
9 3 0 2 3 0 2 3 2 0
10 3 0 3 0 3 1 3 3 0 0
14 3 3 1 3 3 0 3 0 1 1 3 0 3 0
6 3 3 1 0 1 2
2 3 3
10 3 0 3 0 3 1 2 0 0 3
3 3 0 3
6 3 1 1 3 3 0
10 3 0 3 1 0 1 3 3 0 3
2 3 3
4 3 0 3 0
9 3 3 1 0 3 0 1 3 0
3 3 0 3
7 3 0 3 0 3 0 3
4 3 3 1 1
11 3 3 2 1 1 2 1 1 2 0 1
1 3
4 3 3 1 1
2 3 3
2 3 3
7 3 0 3 0 3 1 3
2 3 3
2 3 0
7 3 0 1 3 3 3 0
6 3 3 1 3 3 3
23 3 3 1 1 1 1 3 0 1 0 2 0 1 2 3 0 2 0 3 3 0 1 3
2 3 3
18 3 1 3 0 2 1 3 2 1 1 3 3 0 2 3 0 3 0
6 3 2 0 3 1 3
9 3 3 1 2 3 1 2 0 3
12 3 3 0 0 0 1 0 2 3 0 3 3
2 3 3
6 3 0 2 3 0 1
9 3 1 1 3 3 3 1 3 0
7 3 0 1 3 3 0 1
3 3 0 3
2 3 1
2 3 3
9 3 3 0 0 1 3 1 3 3
1 3
12 3 0 2 3 1 1 1 1 3 1 3 0
3 3 3 0
3 3 0 3
16 3 3 1 3 3 1 2 0 3 0 1 1 2 1 1 3
7 3 3 1 3 3 0 3
5 3 3 2 1 3
9 3 0 2 1 3 0 0 3 3
2 3 3
10 3 3 1 3 3 0 3 0 2 1
7 3 0 3 3 3 0 3
1 3
2 3 3
5 3 1 0 0 0
4 3 3 2 3
3 3 0 3
3 3 1 3
3 3 0 1
5 3 0 3 3 0
18 3 0 3 0 2 1 0 2 0 1 0 1 3 3 0 0 2 3
3 3 0 3
5 3 0 3 3 0
3 3 3 0
5 3 0 3 0 2
10 3 1 3 1 1 1 1 1 1 3
2 3 3
27 3 0 3 0 3 0 0 1 2 3 0 0 0 1 1 2 3 0 0 1 3 0 2 0 1 3 3
17 3 0 3 0 0 1 3 3 1 2 2 3 0 3 3 3 3
20 3 0 2 3 0 1 1 2 3 1 2 3 0 3 0 1 3 3 1 3
3 3 3 2
17 3 1 2 0 2 0 3 1 2 0 3 1 3 1 0 3 0
2 3 3
5 3 1 3 1 2
2 3 3
4 3 0 3 0
3 3 0 3
4 3 1 3 0
8 3 3 1 3 3 1 3 3
4 3 0 0 3
7 3 3 0 2 3 2 0
3 3 0 3
4 3 1 0 0
13 3 0 3 1 2 3 0 1 0 2 3 3 1
6 3 0 2 3 3 3
4 3 3 0 0
14 3 0 3 1 2 1 1 1 1 1 1 1 1 0
8 3 0 2 1 3 0 0 0
10 3 1 3 0 2 0 3 0 0 2
2 3 3
3 3 1 0
2 3 3
4 3 1 3 0
8 3 3 0 2 2 0 1 3
3 3 0 3
12 3 0 0 2 3 1 0 0 3 0 2 0
3 3 3 0
1 3
9 3 0 3 0 1 2 2 0 3
3 3 0 1
7 3 0 3 0 1 2 3
6 3 3 2 2 2 3
3 3 0 3
13 3 0 3 0 1 0 1 2 2 3 1 3 3
1 3
7 3 3 0 0 3 3 1
7 3 1 1 3 0 3 3
14 3 1 3 0 0 3 3 3 3 3 1 3 3 2
2 3 0
13 3 3 1 1 3 2 2 0 3 0 1 1 3
3 3 2 1
2 3 3
15 3 3 3 0 0 3 1 3 3 3 0 1 3 3 3
3 3 3 0
20 3 1 1 1 1 1 1 1 1 1 3 1 1 3 0 0 3 3 0 3
9 3 3 0 1 3 0 1 3 1
21 3 3 3 0 3 3 3 0 3 0 1 0 3 3 0 1 3 3 1 2 3
2 3 3
1 3
4 3 1 2 0
8 3 3 0 0 3 3 1 2
12 3 0 3 3 1 3 3 2 0 1 1 3
6 3 0 3 0 1 0
3 3 0 3
5 3 1 3 1 1
3 3 3 0
3 3 0 2
2 3 3
3 3 1 3
12 3 3 0 1 2 0 3 3 1 1 2 1
5 3 3 2 0 3
7 3 0 3 1 3 0 3
2 3 3
2 3 3
6 3 0 3 0 0 1
4 3 1 3 0
28 3 0 3 0 0 2 2 3 2 3 0 1 3 3 0 3 0 1 1 3 2 2 0 3 0 1 3 3
19 3 3 1 3 3 1 3 0 0 1 2 2 0 3 0 2 1 0 1
2 3 3
1 3
2 3 3
7 3 1 1 3 1 0 0
6 3 3 0 2 1 2
21 3 0 3 0 2 3 1 2 0 3 1 2 3 0 1 1 1 2 3 0 0
4 3 3 2 0
16 3 0 3 1 2 2 0 3 1 2 0 1 3 0 0 3
22 3 1 3 1 3 1 3 1 3 3 3 0 2 3 1 1 1 2 1 3 3 2
12 3 0 3 0 1 3 3 1 2 0 3 0
12 3 3 1 3 3 3 1 2 3 0 2 3
10 3 0 3 0 1 1 1 1 1 0
1 3
13 3 0 3 0 1 1 3 3 0 2 3 2 0
14 3 1 1 1 3 3 3 0 2 0 3 0 1 3
3 3 0 3
26 3 3 1 3 3 1 0 2 1 1 2 0 3 0 2 1 3 0 0 1 1 3 0 1 1 0
7 3 3 1 3 3 0 3
5 3 3 0 0 0
4 3 0 3 0
25 3 0 3 0 1 2 1 3 2 1 3 1 1 0 3 3 0 3 0 0 3 3 3 3 3
8 3 1 3 1 3 0 0 0
3 3 3 3
18 3 0 3 0 1 3 3 1 2 1 2 0 3 0 3 0 2 0
4 3 0 3 3
4 3 3 1 2
2 3 3
10 3 3 1 3 3 1 3 3 1 1
4 3 0 2 3
1 3
10 3 0 1 2 1 1 2 1 3 0
7 3 3 3 1 3 0 0
25 3 3 0 1 3 1 1 2 1 1 1 1 1 2 3 1 3 3 0 3 0 1 0 3 0
13 3 1 1 3 3 0 1 3 3 1 2 1 3
9 3 0 2 3 0 1 2 3 2
10 3 3 0 0 1 3 0 0 1 3
11 3 0 3 0 3 0 1 2 0 1 1
9 3 3 0 2 0 3 1 2 3
3 3 3 2
5 3 1 2 0 0
1 3
11 3 1 3 3 0 3 0 1 3 3 3
9 3 0 3 0 3 0 2 0 3
4 3 3 1 0
9 3 1 3 0 0 1 1 3 0
3 3 1 3
3 3 1 0
5 3 3 1 3 1
22 3 3 0 2 3 1 3 3 0 1 0 1 3 3 1 2 1 2 3 1 3 3
4 3 0 3 3
23 3 0 3 1 2 1 1 1 1 1 1 2 3 1 0 0 1 2 2 3 3 2 0
7 3 2 0 2 3 0 2
6 3 3 1 3 3 0
3 3 0 3
7 3 1 1 1 3 0 1
6 3 0 3 0 2 3
5 3 0 1 1 1
3 3 1 3
3 3 3 0
4 3 0 2 3
7 3 0 3 1 1 3 0
15 3 0 3 0 1 3 3 0 0 2 1 1 2 0 1
23 3 0 3 3 3 1 0 0 1 3 3 3 0 1 1 3 3 1 1 1 2 0 3
6 3 1 2 1 3 0
2 3 3
12 3 0 0 2 0 1 3 0 2 3 2 3
11 3 3 1 3 3 0 1 3 3 3 0
5 3 3 0 0 3
3 3 1 3
6 3 3 0 0 0 1
10 3 1 3 0 2 0 3 3 2 0
3 3 3 2
6 3 3 1 3 3 3
2 3 3
2 3 3
2 3 2
6 3 0 3 3 0 1
2 3 3
37 3 3 1 3 3 0 2 1 1 1 1 3 0 1 1 1 2 0 3 1 3 0 3 0 1 3 3 0 3 0 3 1 2 2 0 1 0
3 3 3 0
26 3 3 1 3 3 0 1 1 1 1 3 2 0 2 0 0 3 1 3 0 3 0 1 3 3 3
13 3 1 3 0 1 0 1 2 3 1 1 1 1
7 3 3 1 3 1 1 3
17 3 1 0 1 1 3 0 2 0 0 2 3 1 3 3 1 0
8 3 3 3 1 3 0 3 3
2 3 3
10 3 0 3 1 2 0 2 0 1 3
3 3 0 1
19 3 3 1 3 3 0 0 3 0 1 2 1 2 3 1 3 3 3 2
9 3 3 1 3 3 1 3 3 2
11 3 3 1 3 3 1 3 0 2 2 2
6 3 3 3 0 0 0
3 3 3 0
6 3 0 3 3 0 2
6 3 3 0 1 1 1
23 3 0 2 2 1 1 2 0 3 0 3 0 3 1 3 3 1 3 3 0 3 0 2
6 3 1 0 1 3 0
2 3 3
4 3 0 3 3
1 3
14 3 3 0 0 0 2 0 3 1 3 0 3 1 3
3 3 0 3
1 3
2 3 3
22 3 1 3 0 1 3 2 2 3 1 3 3 1 2 0 3 1 3 3 0 0 2
2 3 3
17 3 3 1 3 3 3 0 0 0 3 3 3 3 0 2 1 2
1 3
6 3 3 2 0 0 0
2 3 3
1 3
8 3 3 1 3 3 0 3 0
8 3 3 1 3 3 1 2 3
3 3 3 0
8 3 3 3 3 3 0 3 0
12 3 3 0 2 0 3 1 2 1 0 2 3
8 3 0 3 0 1 3 3 0
3 3 3 1
20 3 1 3 0 2 1 1 3 3 0 1 2 3 1 2 1 3 1 0 0
6 3 3 1 3 3 3
9 3 2 0 0 1 3 0 0 3
14 3 3 1 2 1 1 1 1 1 1 1 1 1 0
8 3 1 3 1 3 3 0 3
13 3 1 2 0 3 1 3 0 3 0 2 0 3
3 3 1 3
4 3 0 3 3
2 3 3
5 3 0 3 2 1
3 3 3 2
2 3 0
10 3 0 3 0 2 3 0 2 0 2
4 3 1 3 0
3 3 1 3
1 3
3 3 1 3
14 3 3 1 3 2 3 3 0 1 1 1 1 2 3
6 3 3 0 1 1 0
4 3 3 3 0
8 3 0 3 1 0 1 3 3
1 3
6 3 0 3 1 0 2
3 3 1 3
5 3 1 2 0 2
2 3 3
3 3 1 3
3 3 3 0
3 3 0 3
2 3 2
5 3 0 2 3 1
5 3 1 1 2 3
14 3 0 3 3 3 0 2 3 1 3 3 0 3 0
3 3 1 2
6 3 1 1 3 0 2
3 3 1 3
2 3 3
5 3 1 1 3 0
12 3 3 0 2 0 3 0 1 1 1 3 0
13 3 0 3 0 1 3 3 3 1 3 3 3 2
9 3 0 3 0 3 0 1 2 3
11 3 3 1 2 1 1 1 1 1 1 1
6 3 0 2 3 0 0
2 3 3
8 3 1 3 0 2 1 2 0
14 3 3 1 3 2 2 0 1 3 0 0 1 3 0
3 3 1 2
3 3 3 0
1 3
1 3
16 3 1 1 3 1 3 0 1 2 3 2 1 1 2 1 1
4 3 3 1 3
12 3 0 3 1 0 1 0 1 3 3 0 0
3 3 1 3
4 3 0 2 3
12 3 3 1 3 3 0 3 1 3 3 2 0
17 3 0 3 0 1 3 3 3 1 3 3 0 3 1 3 1 3
6 3 0 3 1 3 3
3 3 0 1
3 3 3 2
10 3 3 2 1 3 3 3 1 1 2
16 3 0 3 1 2 2 3 2 0 2 1 1 3 2 0 3
3 3 0 3
5 3 2 0 3 0
21 3 0 2 3 0 2 2 0 0 3 0 0 1 3 0 0 3 0 3 2 1
3 3 3 0
24 3 0 3 1 2 1 1 2 3 1 3 3 1 1 3 3 0 3 0 3 1 2 1 3
3 3 3 0
5 3 1 3 1 1
2 3 3
2 3 3
4 3 0 3 0
3 3 3 0
9 3 3 1 3 3 1 3 3 2
5 3 0 3 3 1
3 3 3 0
3 3 3 1
7 3 0 3 3 0 2 3
3 3 1 2
13 3 0 3 0 1 3 3 3 0 2 1 1 3
5 3 0 3 1 2
6 3 3 3 1 3 3
4 3 0 3 3
4 3 3 1 0
4 3 2 0 2
3 3 1 3
8 3 0 3 3 3 0 2 0
5 3 1 3 0 1
28 3 1 1 3 1 3 3 0 1 3 3 0 3 0 1 3 3 0 1 3 3 0 3 0 3 1 2 3
3 3 3 0
3 3 1 3
7 3 1 1 1 3 3 0
15 3 0 3 1 0 1 2 1 1 1 1 2 0 2 3
11 3 0 3 0 2 3 3 1 3 3 3
10 3 3 1 3 3 3 1 3 1 2
5 3 1 3 0 1
4 3 0 0 0
4 3 1 1 3
4 3 0 3 0
2 3 3
6 3 3 0 2 0 3
11 3 3 0 3 3 0 3 0 2 0 3
4 3 0 2 3
4 3 3 0 3
4 3 3 0 2
6 3 0 3 3 2 1
4 3 0 3 3
5 3 0 3 1 3
22 3 1 2 0 2 3 1 3 0 1 2 0 3 0 0 3 1 3 3 1 3 1
9 3 3 2 1 3 0 2 2 3
3 3 1 3
4 3 0 3 3
3 3 3 2
9 3 3 3 1 3 0 2 1 2
3 3 3 2
7 3 0 3 0 2 0 3
7 3 3 0 2 0 1 0
11 3 3 2 0 3 0 0 3 0 2 0
2 3 2
10 3 3 1 2 0 0 1 3 3 3
3 3 0 3
5 3 3 3 2 1
1 3
4 3 3 2 0
7 3 0 3 0 2 0 0
8 3 0 3 3 1 3 3 3
5 3 2 0 3 0
20 3 3 3 3 0 1 2 1 1 2 1 1 3 1 3 3 1 0 3 3
2 3 1
3 3 0 3
3 3 0 3
3 3 3 0
2 3 0
2 3 3
6 3 0 3 0 2 0
3 3 3 2
2 3 3
1 3
2 3 3
7 3 1 2 0 0 1 3
3 3 0 3
19 3 0 3 1 3 0 3 0 1 3 3 3 1 1 1 3 1 3 0
17 3 0 3 1 2 2 0 3 3 1 3 3 3 0 3 3 0
1 3
24 3 0 1 3 3 3 0 2 1 3 0 2 0 3 1 0 2 0 0 2 3 1 3 2
2 3 1
14 3 3 1 3 3 3 0 0 1 1 1 1 3 0
3 3 0 3
5 3 1 3 0 2
11 3 0 2 3 0 2 1 1 1 3 0
5 3 0 2 0 1
2 3 3
5 3 0 3 1 3
3 3 1 3
18 3 0 3 0 1 0 1 1 3 3 2 0 0 2 1 1 3 0
25 3 1 3 1 0 1 1 1 2 0 2 3 0 1 1 1 2 0 3 0 1 3 3 0 3
4 3 0 3 3
6 3 0 1 1 1 3
3 3 0 3
2 3 3
9 3 0 3 1 0 2 1 1 0
9 3 3 0 2 0 2 2 2 3
2 3 3
2 3 3
6 3 3 0 2 3 3
4 3 1 3 0
1 3
4 3 1 3 2
12 3 3 2 0 1 0 2 0 0 2 3 3
10 3 0 3 0 1 3 3 3 0 2
4 3 1 3 0
2 3 3
7 3 3 3 3 1 3 0
19 3 0 3 0 0 3 1 3 3 0 1 3 2 0 3 0 1 1 3
10 3 0 3 1 3 0 0 2 3 0
2 3 3
3 3 0 3
4 3 3 1 3
12 3 0 3 0 1 2 2 0 3 0 3 3
6 3 0 3 0 1 2
3 3 3 2
3 3 0 1
3 3 3 0
4 3 3 0 3
1 3
14 3 3 2 3 2 0 3 1 3 3 0 1 3 3
22 3 0 1 0 1 3 1 3 3 0 1 1 0 3 3 3 3 3 3 0 2 1
4 3 0 2 3
13 3 0 2 3 0 1 3 0 1 3 3 0 2
9 3 3 1 3 3 1 0 2 3
11 3 0 3 0 2 1 0 1 3 3 3
2 3 3
10 3 3 0 2 1 3 3 1 1 3
3 3 0 3
9 3 3 1 1 1 1 1 1 3
2 3 3
5 3 2 0 3 0
2 3 1
5 3 1 3 0 2
7 3 3 2 0 0 3 3
17 3 0 3 1 2 1 1 1 3 0 0 1 3 0 2 0 3
1 3
1 3
3 3 1 3
3 3 1 3
5 3 0 2 3 0
3 3 3 0
10 3 0 3 0 1 2 0 3 3 3
26 3 0 3 1 2 1 1 1 1 1 2 3 1 3 3 1 0 3 3 0 1 3 1 2 0 3
9 3 0 3 0 2 3 0 2 0
4 3 2 0 3
7 3 2 0 3 0 0 0
2 3 3
17 3 0 3 3 1 3 3 1 2 1 1 1 1 1 2 0 1
7 3 3 0 0 1 3 0
15 3 0 3 3 2 0 2 0 3 0 1 3 3 0 3
3 3 0 1
10 3 3 1 2 1 1 1 3 1 1
11 3 0 3 3 1 3 3 3 1 3 0
3 3 3 0
8 3 3 2 3 1 3 3 0
1 3
2 3 3
3 3 0 3
2 3 3
5 3 0 3 0 0
5 3 3 1 2 3
8 3 0 3 1 3 3 0 0
35 3 3 0 1 0 1 3 0 3 2 0 1 2 1 2 3 1 2 3 0 3 1 2 1 1 3 0 1 3 3 0 2 2 1 3
3 3 0 0
2 3 3
18 3 0 3 0 1 3 3 3 0 2 3 1 1 0 1 1 1 3
11 3 0 2 3 0 2 0 3 0 3 3
1 3
5 3 0 3 1 2
9 3 0 3 1 2 1 1 1 3
6 3 3 3 1 3 3
5 3 0 3 1 3
1 3
7 3 1 3 0 0 1 3
13 3 0 3 0 3 0 1 2 1 1 1 1 0
1 3
8 3 0 3 1 2 0 1 3
2 3 3
17 3 1 3 0 1 2 0 2 3 1 1 1 1 1 1 1 2
10 3 3 0 1 3 2 2 0 2 3
8 3 3 0 3 3 2 0 0
2 3 3
4 3 3 0 1
5 3 1 1 1 3
14 3 3 0 2 2 0 3 0 2 1 3 1 3 3
5 3 1 3 0 2
3 3 3 2
8 3 1 3 0 1 1 1 0
8 3 0 3 0 3 3 0 2
3 3 3 0
7 3 3 1 2 3 3 0
11 3 3 1 3 1 3 1 3 3 0 3
2 3 3
13 3 1 3 1 3 3 1 2 3 0 1 1 1
9 3 3 1 3 3 0 3 3 1
12 3 3 0 1 2 0 3 1 3 2 0 0
12 3 0 3 0 1 3 3 0 1 2 0 3
7 3 3 1 3 3 1 3
5 3 0 1 3 3
7 3 1 2 0 0 1 3
2 3 3
1 3
27 3 0 3 3 0 1 1 1 1 2 0 3 1 2 0 1 3 0 1 3 0 3 2 1 3 2 3
10 3 0 3 3 1 3 1 1 1 0
9 3 3 0 0 0 3 3 1 0
10 3 0 3 0 3 0 1 3 2 0
1 3
7 3 3 1 1 3 3 3
15 3 3 0 0 3 3 3 3 3 0 1 3 3 1 3
1 3
21 3 0 3 1 0 1 2 3 1 0 0 1 3 3 3 0 3 1 3 0 3
8 3 0 2 3 3 3 3 3
2 3 1
7 3 3 0 2 3 1 3
3 3 1 0
6 3 3 1 3 3 3
1 3
14 3 3 0 1 2 0 3 0 2 3 0 1 0 2
15 3 0 1 1 1 1 2 3 0 0 2 3 2 0 3
2 3 1
2 3 3
19 3 1 3 1 3 3 0 3 3 0 0 0 3 3 3 0 0 2 3
6 3 0 0 2 1 3
16 3 3 1 3 3 0 3 0 1 2 3 3 1 0 3 0
4 3 0 2 3
3 3 3 0
6 3 1 1 3 0 0
39 3 0 3 0 3 0 1 0 1 3 3 3 1 3 3 0 2 0 1 3 3 1 3 0 2 0 1 3 3 0 3 0 1 2 1 2 3 0 2
5 3 3 0 0 0
8 3 0 3 1 3 1 1 3
15 3 3 2 0 2 1 3 2 0 0 3 3 0 3 0
5 3 0 3 1 3
3 3 0 3
10 3 0 3 0 1 2 1 3 3 3
6 3 0 3 0 0 3
9 3 3 0 1 1 3 1 2 3
8 3 3 0 1 2 1 1 3
2 3 3
16 3 0 2 3 0 2 2 0 1 3 0 1 3 2 1 3
5 3 0 3 3 0
2 3 0
1 3
2 3 3
16 3 3 0 0 0 3 3 3 0 3 1 2 2 1 3 0
14 3 3 0 0 3 3 0 2 3 1 0 1 3 0
1 3
12 3 0 3 0 1 0 0 1 1 2 0 3
5 3 3 1 1 0
10 3 0 3 0 2 3 1 3 3 3
22 3 3 0 2 1 2 3 1 3 3 0 1 2 0 1 1 3 1 2 3 0 3
12 3 0 3 0 1 0 1 2 1 1 0 2
2 3 3
3 3 0 3
13 3 3 1 2 1 0 0 0 3 0 1 2 0
11 3 3 0 2 0 3 0 2 2 2 3
12 3 1 3 0 2 1 2 0 1 0 1 1
10 3 0 3 0 3 1 2 3 0 0
17 3 1 3 0 3 3 3 0 3 0 2 0 0 1 3 3 3
9 3 1 1 1 3 1 1 1 2
1 3
13 3 3 2 3 0 2 3 3 2 3 3 0 0
9 3 0 3 0 3 1 3 1 3
8 3 3 0 2 1 3 3 2
9 3 1 0 1 1 3 0 0 3
3 3 3 2
8 3 3 0 2 0 3 1 1
2 3 3
6 3 1 2 0 0 0
5 3 2 0 3 1
6 3 0 3 1 2 3
3 3 0 3
12 3 3 1 3 3 1 3 0 2 1 3 0
17 3 0 3 0 2 0 0 1 0 2 3 1 2 3 0 2 0
11 3 1 1 3 3 3 1 3 3 0 2
6 3 1 1 3 0 0
12 3 3 1 3 3 0 2 1 0 1 3 3
16 3 0 3 1 2 1 2 0 3 1 0 2 0 3 1 3
5 3 0 3 0 2
17 3 1 1 3 1 1 3 0 1 1 3 2 0 3 1 3 3
3 3 0 3
5 3 3 1 3 2
19 3 1 2 0 1 1 2 3 1 3 3 0 3 1 0 1 2 3 0
6 3 1 0 1 3 0
5 3 0 3 3 0
6 3 3 1 1 0 0
6 3 1 3 0 2 1
3 3 1 3
10 3 0 3 1 2 2 0 3 0 3
2 3 3
2 3 3
7 3 0 0 2 3 0 0
8 3 0 2 3 0 2 0 3
3 3 1 3
3 3 1 3
4 3 3 0 2
5 3 3 1 3 3
12 3 0 3 0 1 0 2 0 0 1 0 0
1 3
14 3 0 3 0 1 2 3 3 3 0 0 1 1 3
2 3 3
7 3 0 3 1 2 0 3
3 3 0 1
3 3 1 2
2 3 3
13 3 3 0 1 1 2 0 3 1 0 1 0 2
2 3 0
5 3 1 3 0 1
3 3 3 0
16 3 0 3 3 1 3 3 1 0 1 2 3 0 0 1 3
5 3 0 3 3 0
16 3 0 1 2 0 0 3 0 0 1 3 0 2 2 0 3
4 3 0 3 3
4 3 3 0 2
4 3 0 2 3
1 3
9 3 3 1 3 2 0 1 1 3
3 3 3 0
4 3 3 0 1
25 3 0 3 0 1 3 3 0 1 3 3 3 1 3 0 3 3 3 3 3 2 1 3 2 0
1 3
1 3
1 3
7 3 0 3 0 1 3 1
2 3 3
4 3 0 3 0
3 3 1 3
14 3 3 1 3 3 0 3 0 1 2 2 0 3 3
1 3
10 3 3 0 2 2 0 3 0 1 0
18 3 0 3 1 3 0 3 3 1 1 1 3 0 3 3 3 0 3
6 3 3 2 0 0 0
8 3 1 2 0 1 1 0 1
5 3 3 0 0 0
3 3 3 0
5 3 3 1 3 3
4 3 2 0 3
6 3 3 1 3 3 3
10 3 3 0 1 0 0 0 3 0 1
2 3 3
5 3 0 3 0 2
2 3 3
11 3 3 1 2 1 2 0 2 1 1 3
3 3 3 1
4 3 0 2 3
14 3 0 3 0 1 1 3 0 3 3 3 0 3 0
29 3 1 1 3 0 3 1 0 1 3 3 1 2 1 1 1 0 1 3 0 3 0 3 3 0 2 0 2 0
3 3 0 3
6 3 3 1 2 3 3
17 3 0 3 0 3 1 2 0 3 0 0 0 1 3 3 3 3
1 3
13 3 3 2 0 0 0 3 3 0 3 1 0 1
7 3 0 2 3 0 0 0
12 3 0 3 0 2 0 3 1 3 3 0 3
6 3 3 0 1 2 0
3 3 1 2
10 3 0 2 3 0 1 3 3 0 2
1 3
9 3 0 3 2 0 3 1 3 3
16 3 0 3 0 2 3 1 3 0 3 1 2 1 1 3 3
3 3 3 0
13 3 3 1 0 3 1 1 3 3 3 0 0 3
2 3 3
3 3 0 3
13 3 3 1 2 2 0 3 0 0 3 1 2 3
2 3 3
8 3 0 3 0 1 2 0 3
5 3 0 3 1 3
2 3 3
10 3 3 0 1 1 3 1 3 0 0
7 3 3 0 1 1 1 0
9 3 1 3 0 2 1 3 1 3
5 3 0 3 0 3
7 3 0 3 1 2 0 3
3 3 0 3
1 3
4 3 0 1 2
11 3 3 3 3 2 1 1 1 2 3 2
3 3 3 3
12 3 0 3 0 1 1 1 3 0 3 3 3
3 3 3 0
4 3 0 3 3
2 3 1
11 3 0 3 0 3 1 3 3 0 2 1
9 3 0 3 0 3 0 0 0 2
3 3 3 0
2 3 2
8 3 0 3 0 1 2 0 3
6 3 0 3 0 1 2
7 3 0 1 0 2 3 0
2 3 3
7 3 0 3 0 0 2 3
2 3 3
4 3 0 3 0
5 3 3 1 0 3
8 3 0 2 3 0 1 1 0
3 3 3 0
3 3 0 3
11 3 0 1 3 3 0 1 1 3 3 0
3 3 3 0
8 3 0 2 3 0 0 1 3
2 3 0
4 3 0 3 0
3 3 0 3
3 3 0 3
2 3 3
14 3 0 3 1 2 2 0 3 0 1 2 1 1 3
2 3 3
17 3 3 1 3 3 0 1 3 3 1 3 0 1 1 1 1 1
17 3 0 3 0 1 3 3 0 3 0 1 1 1 3 1 1 3
22 3 0 3 1 3 0 3 0 1 1 3 1 3 0 2 1 2 0 1 2 1 3
4 3 3 1 0
10 3 3 0 1 2 0 3 2 0 3
2 3 3
2 3 0
2 3 0
44 3 0 3 0 1 3 3 3 1 3 3 3 0 1 3 1 1 0 1 3 2 2 1 0 3 3 3 3 3 0 3 1 0 2 0 0 1 1 1 1 3 1 3 1
5 3 2 0 3 0
8 3 1 3 0 2 2 0 3
7 3 0 3 3 1 3 3
7 3 0 3 0 1 3 3
11 3 0 2 3 1 3 2 1 1 2 0
7 3 1 2 2 0 3 0
6 3 1 1 3 0 3
19 3 0 3 1 3 0 3 0 1 3 3 3 0 2 3 1 3 3 3
5 3 3 2 3 0
4 3 2 0 3
3 3 1 0
10 3 0 3 0 1 3 2 1 3 3
2 3 3
20 3 0 3 1 3 0 0 1 3 2 0 1 3 3 3 1 3 3 3 0
11 3 1 1 3 1 3 3 1 2 0 3
8 3 0 3 0 3 1 0 2
2 3 0
5 3 3 0 1 1
2 3 0
7 3 3 0 0 1 3 0
5 3 1 3 0 0
2 3 3
1 3
3 3 0 1
5 3 0 3 1 3
1 3
6 3 1 0 3 3 0
9 3 0 3 1 2 0 3 0 2
3 3 0 3
1 3
3 3 1 3
8 3 0 3 3 0 2 3 1
19 3 0 3 0 0 2 0 3 0 1 3 3 3 1 2 2 0 0 2
10 3 0 3 0 1 3 3 1 1 3
30 3 3 0 2 0 3 0 1 1 3 3 0 1 3 3 3 0 2 0 3 0 1 2 3 3 0 2 0 3 3
4 3 3 1 3
2 3 0
4 3 1 3 0
4 3 3 0 1
5 3 0 0 2 3
8 3 3 0 3 1 1 3 3
5 3 1 2 1 2
5 3 3 0 0 0
5 3 3 1 0 0
12 3 1 3 1 3 3 0 2 2 2 3 0
3 3 1 3
14 3 0 3 0 1 2 1 1 1 2 3 0 0 2
13 3 0 3 0 3 0 1 3 3 3 2 3 3
5 3 0 3 1 3
2 3 0
2 3 3
5 3 1 2 1 3
7 3 0 3 1 3 2 1
8 3 0 2 3 0 1 2 3
1 3
13 3 3 1 3 3 3 0 1 1 0 3 0 0
3 3 3 0
2 3 3
6 3 3 2 3 0 3
3 3 3 0
15 3 0 3 0 3 0 0 3 1 3 3 0 3 3 0
10 3 2 3 0 1 3 3 1 2 3
5 3 3 1 3 3
5 3 0 2 0 3
12 3 0 3 1 3 0 3 1 2 0 3 0
6 3 3 1 3 3 0
2 3 3
4 3 0 3 0
3 3 0 3
1 3
2 3 3
3 3 0 2
19 3 3 1 1 0 2 3 3 1 3 3 1 3 3 3 0 1 2 3
16 3 0 1 2 3 3 1 3 1 3 1 3 3 1 1 1
6 3 3 1 3 3 3
13 3 0 3 1 2 3 0 2 1 0 3 3 3
5 3 0 3 0 3
2 3 3
3 3 0 3
12 3 0 3 0 1 3 3 0 3 3 0 2
13 3 3 1 3 3 3 0 1 3 2 0 1 3
8 3 3 0 2 0 3 3 0
8 3 3 1 2 3 0 3 0
3 3 0 3
2 3 3
2 3 3
4 3 0 3 3
9 3 3 1 3 3 0 3 0 3
9 3 0 3 0 3 0 2 0 0
4 3 0 2 3
8 3 3 0 0 1 1 3 0
5 3 1 3 0 0
3 3 0 3
2 3 3
6 3 0 3 0 3 0
4 3 2 0 1
10 3 1 0 0 0 1 1 3 3 0
3 3 1 3
19 3 1 3 0 2 0 2 2 2 0 3 0 1 2 3 0 2 1 2
9 3 0 3 1 0 2 1 3 3
13 3 0 3 1 1 3 3 0 2 3 2 0 3
4 3 1 3 0
10 3 1 1 3 1 3 3 3 0 3
3 3 1 3
5 3 1 1 3 3
5 3 1 3 0 0
8 3 0 2 3 0 1 0 1
12 3 3 0 3 0 3 0 1 3 3 0 3
2 3 3
3 3 0 3
2 3 3
12 3 0 3 0 0 3 1 2 2 0 3 3
13 3 3 0 2 0 1 2 3 1 1 1 3 0
3 3 0 3
2 3 3
1 3
6 3 0 3 0 1 3
2 3 3
12 3 3 0 1 1 2 3 1 3 3 1 3
5 3 0 3 0 1
1 3
5 3 3 1 0 0
4 3 3 0 3
10 3 1 0 0 3 3 3 3 1 0
2 3 3
3 3 0 1
16 3 3 0 2 2 0 3 1 3 2 1 1 2 0 3 3
18 3 0 3 0 1 3 3 3 0 2 0 3 1 3 1 3 0 0
17 3 0 3 1 2 0 3 0 1 1 1 1 3 1 3 3 3
2 3 3
2 3 1
6 3 0 3 0 3 0
4 3 3 0 2
9 3 3 1 0 0 2 0 3 3
13 3 3 1 3 3 1 1 3 3 0 2 1 3
9 3 1 3 1 3 3 0 1 2
21 3 0 3 0 2 3 0 1 0 3 3 3 3 1 2 0 3 0 2 0 3
3 3 1 3
3 3 0 3
2 3 3
12 3 0 3 0 1 1 1 1 1 1 1 1
5 3 3 0 2 3
1 3
13 3 0 3 0 1 1 3 2 3 1 2 3 0
2 3 3
2 3 3
3 3 0 3
6 3 0 3 0 0 3
8 3 0 3 0 2 3 1 2
8 3 3 1 3 3 1 2 3
22 3 0 3 0 2 3 1 1 3 0 2 3 1 1 0 1 3 1 0 1 3 3
5 3 3 0 1 0
5 3 3 1 3 3
20 3 0 1 2 2 0 3 1 3 3 0 0 2 1 1 3 1 3 3 3
15 3 3 1 3 1 2 1 0 3 3 1 2 1 1 3
31 3 0 3 1 3 0 3 0 1 3 1 1 1 1 3 2 1 1 3 3 0 0 1 0 0 3 3 3 0 2 3
5 3 0 3 0 3
6 3 1 3 0 1 1
7 3 0 3 1 2 1 3
3 3 1 3
3 3 0 3
13 3 0 3 1 3 0 0 3 3 1 0 2 0
5 3 0 3 0 3
17 3 3 1 1 3 0 1 3 3 3 1 1 3 3 1 2 3
17 3 3 1 3 3 1 1 1 1 3 0 2 1 3 2 0 2
10 3 3 1 3 2 0 3 3 3 2
4 3 3 2 2
10 3 0 3 0 1 0 0 3 3 3
2 3 3
6 3 0 3 0 1 2
2 3 3
10 3 0 3 1 2 1 1 1 2 3
10 3 0 3 1 2 1 2 1 1 2
6 3 3 0 2 0 1
3 3 3 3
2 3 3
3 3 0 3
22 3 0 3 3 0 3 3 0 3 0 0 3 0 2 1 0 1 2 1 1 0 0
5 3 3 1 0 0
11 3 3 0 1 1 3 3 3 3 3 1
16 3 0 2 1 0 0 3 1 0 1 3 3 3 1 0 0
9 3 3 0 2 1 0 3 3 3
6 3 0 3 1 0 2
6 3 2 0 3 0 1
3 3 0 3
8 3 0 3 0 1 1 3 3
33 3 0 3 1 0 1 3 3 3 0 0 2 1 3 0 1 2 0 3 0 1 3 3 0 1 1 1 1 1 2 3 1 2
14 3 1 3 0 2 0 3 1 3 3 2 1 1 1
2 3 3
3 3 1 3
1 3
9 3 3 0 1 1 3 0 1 3
2 3 3
3 3 3 3
6 3 0 3 0 3 0
4 3 0 2 3
4 3 3 0 0
19 3 3 1 3 3 1 3 0 3 1 0 2 3 2 0 3 0 0 0
2 3 3
13 3 0 1 0 1 0 3 1 0 3 0 1 0
3 3 3 0
10 3 1 1 3 3 0 1 2 3 1
6 3 3 3 2 0 0
1 3
10 3 0 3 1 3 0 3 1 3 1
1 3
10 3 1 3 0 2 3 1 3 3 3
7 3 0 3 1 3 3 3
4 3 0 2 3
2 3 0
10 3 0 3 1 2 1 1 2 0 3
3 3 3 0
15 3 1 3 0 3 3 3 0 3 0 1 0 1 0 2
11 3 1 0 3 3 0 3 1 0 1 3
3 3 3 0
2 3 3
13 3 0 3 0 3 1 2 0 3 0 2 0 3
2 3 3
5 3 1 3 0 0
8 3 0 2 3 0 0 1 3
6 3 0 2 1 3 0
2 3 0
12 3 0 3 0 1 2 3 0 2 2 0 3
2 3 3
13 3 0 3 1 2 3 0 2 0 1 2 1 3
3 3 0 3
6 3 3 1 2 1 1
4 3 0 3 3
4 3 1 3 0
7 3 3 1 3 0 3 0
8 3 3 2 1 3 3 3 0
4 3 3 1 3
5 3 0 3 0 3
6 3 0 1 2 1 0
1 3
15 3 0 1 1 1 1 2 1 1 3 1 0 1 3 3
4 3 3 0 0
11 3 3 1 3 3 0 3 1 0 1 0
15 3 1 3 0 2 3 1 3 3 1 2 2 1 1 0
7 3 1 3 0 2 0 3
1 3
22 3 0 3 1 1 3 3 0 3 0 2 3 0 1 3 3 3 1 3 3 0 0
2 3 3
1 3
3 3 3 2
11 3 1 1 0 0 2 2 0 1 3 0
6 3 3 0 1 2 0
9 3 0 3 0 3 0 2 3 0
27 3 3 1 0 3 3 0 0 3 0 2 3 0 1 0 3 1 3 3 0 2 3 3 1 1 1 3
6 3 1 3 0 2 3
1 3
6 3 3 0 0 3 0
2 3 3
16 3 0 3 1 0 1 2 2 0 3 1 2 1 2 0 3
6 3 3 1 3 3 0
11 3 3 0 1 1 1 2 0 3 3 3
6 3 3 0 2 1 2
2 3 3
5 3 3 0 0 0
8 3 1 2 1 0 3 3 3
2 3 3
3 3 0 3
8 3 0 3 1 2 0 3 0
3 3 0 3
11 3 1 3 0 1 2 3 0 2 3 2
2 3 3
4 3 0 3 3
2 3 0
29 3 3 0 2 3 1 3 3 3 1 3 3 3 1 3 0 2 1 1 3 1 3 3 0 3 2 0 3 0
5 3 1 1 3 3
6 3 0 3 1 2 1
24 3 1 1 1 1 1 3 3 0 1 3 3 3 1 3 0 3 0 3 0 3 0 0 3
4 3 3 2 3
1 3
3 3 0 2
10 3 0 3 2 0 3 0 2 1 3
4 3 0 2 3
5 3 0 3 1 3
26 3 1 1 3 3 0 1 0 1 2 1 1 2 0 3 1 2 3 0 2 1 1 3 3 0 3
1 3
3 3 1 2
7 3 0 3 0 2 3 1
5 3 0 3 1 3
3 3 1 3
33 3 3 2 0 3 0 1 1 3 2 3 0 2 0 3 1 0 1 3 3 0 0 3 0 1 1 3 2 1 1 3 1 0
5 3 0 3 3 2
4 3 3 0 2
1 3
7 3 0 2 1 3 0 0
11 3 3 0 2 0 3 3 1 2 0 3
2 3 3
9 3 0 3 0 1 1 3 3 3
5 3 3 1 3 3
18 3 0 3 0 1 3 1 3 0 0 3 3 0 1 2 0 1 3
6 3 3 0 2 0 3
2 3 1
3 3 1 3
8 3 0 2 2 2 3 0 0
3 3 3 2
4 3 3 3 0
4 3 1 3 3
16 3 0 3 0 2 3 0 3 0 2 1 2 0 1 2 0
8 3 1 3 0 0 1 1 3
2 3 3
6 3 3 0 0 1 3
14 3 1 3 0 1 1 1 1 2 0 2 3 0 0
2 3 0
8 3 0 3 0 1 2 3 0
6 3 0 3 0 2 3
1 3
5 3 3 0 1 3
2 3 3
19 3 0 3 0 1 3 3 0 3 1 3 3 1 3 3 3 1 3 3
5 3 3 1 0 3
4 3 1 1 3
17 3 1 0 3 3 1 3 0 0 0 3 3 3 3 1 3 3
3 3 0 3
1 3
24 3 3 0 0 1 1 3 1 3 3 3 0 3 2 0 3 3 1 3 3 1 3 0 0
3 3 1 2
7 3 3 0 1 1 3 1
3 3 1 3
13 3 0 3 0 3 1 0 1 3 3 0 2 3
3 3 1 3
5 3 0 3 1 2
1 3
3 3 0 3
2 3 3
3 3 3 0
2 3 0
2 3 3
23 3 0 3 1 3 0 2 0 3 0 1 0 2 1 0 1 3 3 0 1 3 1 3
5 3 0 3 0 3
4 3 0 3 3
8 3 0 2 3 0 1 2 3
3 3 0 3
7 3 3 1 2 3 1 3
3 3 1 3
5 3 0 3 0 2
10 3 1 3 0 1 1 1 1 1 0
11 3 0 1 2 2 0 3 0 2 0 0
5 3 0 3 0 3
3 3 0 3
3 3 0 3
16 3 0 2 1 1 3 0 1 3 1 0 1 3 0 1 3
12 3 1 3 0 2 1 1 3 3 0 3 0
4 3 1 3 0
2 3 3
6 3 0 2 3 3 0
7 3 0 3 3 1 0 0
9 3 0 3 0 1 3 3 2 1
17 3 3 1 3 3 1 2 1 2 0 3 0 1 3 3 0 2
3 3 0 1
3 3 0 3
1 3
6 3 1 3 0 2 3
5 3 2 1 2 3
6 3 0 3 1 3 3
3 3 0 3
11 3 1 3 0 0 1 0 1 3 3 0
2 3 3
6 3 1 3 1 2 1
19 3 2 0 3 0 2 2 0 3 0 0 0 1 1 1 3 1 1 3
8 3 3 2 1 3 3 1 3
6 3 3 3 1 3 3
11 3 0 3 0 3 3 1 3 3 0 1
4 3 3 0 0
3 3 0 3
23 3 3 0 1 2 3 0 2 0 3 1 2 1 1 1 1 0 1 3 3 3 3 0
6 3 3 0 2 1 0
2 3 1
2 3 3
6 3 0 3 1 2 1
1 3
5 3 0 2 1 3
7 3 3 0 3 3 0 3
4 3 3 2 0
7 3 0 3 0 1 0 0
8 3 0 3 0 1 1 3 3
3 3 0 3
2 3 3
3 3 0 3
3 3 0 3
8 3 3 1 3 0 0 0 3
2 3 0
10 3 3 1 1 0 0 3 0 2 0
4 3 0 3 3
18 3 3 0 0 1 3 0 1 1 0 2 3 1 3 2 3 1 3
19 3 3 0 2 1 1 3 3 0 1 3 3 0 3 1 2 3 0 2
4 3 1 3 0
26 3 0 3 1 3 0 0 1 1 3 0 1 3 0 2 0 3 3 0 0 3 3 2 0 3 3
1 3
18 3 3 0 3 3 0 2 3 0 2 0 3 1 2 3 1 3 3
13 3 3 0 3 3 0 3 0 3 0 2 3 0
6 3 1 3 0 1 0
1 3
3 3 0 3
7 3 3 1 3 3 0 3
3 3 0 3
12 3 0 3 0 1 3 3 0 1 3 3 3
8 3 0 3 1 2 1 3 0
6 3 3 0 1 0 1
1 3
3 3 3 0
3 3 3 2
2 3 0
24 3 3 1 3 3 3 1 3 3 0 0 0 2 1 3 0 2 3 1 3 1 3 0 2
3 3 3 0
5 3 1 3 0 2
9 3 0 3 0 1 2 3 0 0
5 3 0 3 0 2
7 3 0 3 0 1 2 0
2 3 1
29 3 0 3 0 1 3 3 0 2 1 1 2 1 1 2 3 1 3 3 1 2 0 3 0 1 1 3 2 3
4 3 1 0 0
5 3 0 3 0 2
3 3 3 1
5 3 0 3 0 3
2 3 3
12 3 1 3 1 3 3 3 0 1 3 0 0
15 3 3 1 3 3 0 1 2 3 0 0 0 3 3 3
16 3 0 3 1 3 0 3 0 1 0 2 3 1 0 2 3
4 3 1 1 3
6 3 1 3 3 1 3
7 3 2 0 2 0 0 3
9 3 3 3 3 1 3 3 1 3
5 3 1 3 0 1
2 3 3
7 3 3 0 0 3 1 0
17 3 3 1 3 3 3 0 3 3 0 1 1 1 3 1 1 0
3 3 1 3
4 3 0 3 0
2 3 0
9 3 3 0 2 0 3 1 2 3
2 3 3
18 3 0 3 0 1 2 3 0 0 1 3 3 0 1 1 0 0 1
3 3 0 3
2 3 3
3 3 3 3
2 3 3
9 3 3 1 3 3 1 1 1 1
10 3 0 3 1 2 0 1 1 1 3
5 3 0 2 1 3
6 3 0 2 1 3 0
7 3 0 3 0 1 1 0
7 3 0 2 3 2 0 3
7 3 0 3 0 1 0 0
12 3 1 1 3 0 3 1 2 2 0 3 1
2 3 3
8 3 1 2 0 0 1 1 3
7 3 1 3 2 1 3 3
5 3 0 3 1 3
1 3
2 3 3
3 3 0 3
6 3 1 1 3 1 3
3 3 0 1
4 3 3 2 0
2 3 3
2 3 3
2 3 3
23 3 0 3 1 2 0 3 0 2 1 3 0 0 0 3 3 3 3 1 2 1 1 0
9 3 1 3 1 3 3 0 2 3
18 3 1 3 1 1 1 1 3 3 2 1 2 0 2 3 1 3 3
10 3 0 3 1 2 1 1 2 1 3
2 3 3
10 3 0 3 3 1 3 3 1 2 3
11 3 0 3 1 2 1 3 2 0 0 3
1 3
27 3 0 3 1 2 1 2 3 1 3 3 0 1 1 3 0 3 1 0 2 2 3 1 2 3 0 0
7 3 3 2 0 2 0 3
12 3 1 3 0 0 0 1 1 2 2 3 2
3 3 1 2
3 3 3 0
13 3 0 3 1 0 1 0 1 3 3 0 3 0
11 3 0 3 1 2 0 3 3 1 3 0
2 3 3
8 3 3 2 0 1 2 0 3
8 3 3 2 1 0 3 3 3
9 3 1 3 0 0 1 3 0 0
8 3 0 3 1 3 0 3 0
37 3 3 0 3 3 0 3 0 1 2 1 1 3 3 3 0 0 0 0 0 3 3 1 1 3 0 3 3 3 0 1 3 3 1 3 0 3
4 3 0 3 1
4 3 3 0 0
3 3 3 0
21 3 0 3 0 1 3 3 3 1 1 1 1 1 1 1 1 1 2 3 2 0
3 3 3 1
8 3 3 1 3 1 1 3 0
5 3 3 0 0 3
2 3 2
5 3 0 2 1 3
3 3 3 0
5 3 2 0 0 3
5 3 0 3 0 3
4 3 1 1 3
1 3
9 3 3 0 3 3 3 0 3 0
7 3 3 1 3 3 1 0
32 3 3 1 3 3 1 3 1 3 3 3 0 0 0 3 1 3 2 0 1 3 0 2 3 0 3 3 0 3 3 0 0
10 3 3 1 3 3 1 2 1 3 0
5 3 0 2 3 1
3 3 3 2
2 3 3
14 3 0 3 1 2 2 0 2 3 1 3 3 0 1
4 3 2 0 3
3 3 1 3
6 3 0 3 1 3 3
6 3 0 3 0 1 2
4 3 3 0 2
2 3 0
3 3 3 0
7 3 3 0 3 3 0 3
15 3 0 3 0 3 0 1 3 3 0 3 1 2 0 3
2 3 3
2 3 3
3 3 1 2
12 3 3 0 3 3 1 1 3 0 1 1 3
9 3 0 3 1 2 2 0 2 3
2 3 0
2 3 3
7 3 0 3 0 1 2 1
9 3 0 3 0 1 3 3 1 3
11 3 0 3 0 3 1 2 1 3 0 0
11 3 0 1 3 3 0 1 3 3 1 3
8 3 3 1 3 3 0 2 3
2 3 3
1 3
16 3 1 0 0 1 3 3 0 1 1 2 0 3 0 3 0
6 3 3 0 2 0 1
15 3 3 1 3 3 3 0 3 0 3 1 3 1 3 1
14 3 0 3 1 2 3 0 2 1 0 1 1 3 0
2 3 3
6 3 2 2 3 1 3
5 3 1 3 0 2
7 3 0 3 1 3 3 0
2 3 2
8 3 3 0 0 0 2 0 3
13 3 0 3 0 3 0 1 3 3 0 2 0 3
11 3 3 1 3 3 0 1 3 3 0 2
3 3 0 3
3 3 0 2
10 3 3 0 2 3 1 3 3 0 3
3 3 3 2
5 3 1 1 3 0
3 3 0 3
17 3 3 0 2 0 3 1 2 1 1 2 0 3 1 3 1 3
16 3 0 1 3 3 3 0 1 0 2 1 3 2 0 0 3
26 3 0 3 0 3 1 2 2 0 3 1 3 0 0 1 3 0 1 1 1 1 2 3 2 0 2
1 3
2 3 3
2 3 0
10 3 3 0 1 1 2 0 0 2 3
11 3 3 1 3 3 3 0 2 0 3 0
9 3 0 3 1 2 0 0 1 3
5 3 0 2 3 0
11 3 0 3 3 3 0 1 1 1 1 2
10 3 3 0 2 1 3 1 3 0 3
2 3 3
5 3 3 2 1 0
2 3 3
3 3 1 3
4 3 0 1 2
4 3 2 0 3
2 3 3
21 3 0 3 1 2 3 1 2 1 3 3 3 1 3 0 2 3 0 0 3 0
1 3
5 3 0 2 1 3
5 3 0 3 1 3
2 3 3
3 3 1 2
5 3 1 2 0 0
6 3 0 1 3 3 0
4 3 0 3 0
4 3 1 1 3
11 3 0 3 0 1 0 0 0 2 0 3
7 3 0 3 1 2 0 3
7 3 3 0 0 1 1 3
4 3 1 3 0
2 3 3
2 3 3
8 3 3 2 0 1 3 2 1
6 3 0 3 1 3 0
8 3 0 2 0 0 1 2 3
3 3 0 3
9 3 1 1 1 3 1 3 1 3
4 3 3 1 1
2 3 1
15 3 3 1 3 3 3 1 1 3 1 3 0 0 3 0
10 3 0 3 0 1 2 3 0 1 3
5 3 0 3 0 2
6 3 3 0 2 1 2
8 3 3 1 1 1 1 3 0
1 3
9 3 1 2 1 3 3 0 2 3
2 3 3
14 3 0 2 1 3 0 2 0 3 1 3 0 2 2
3 3 1 3
11 3 3 0 2 3 3 0 0 1 3 0
7 3 3 0 0 1 3 0
2 3 3
3 3 0 0
2 3 3
6 3 0 3 1 2 3
4 3 0 3 0
1 3
6 3 0 3 0 1 3
6 3 0 3 0 0 2
6 3 3 1 3 3 1
21 3 1 1 3 1 3 1 3 0 1 1 1 3 2 1 1 3 3 0 2 0
2 3 3
4 3 0 2 2
4 3 3 0 2
11 3 3 2 0 0 1 3 0 0 1 3
5 3 2 0 3 0
13 3 0 3 1 0 1 3 1 2 3 2 0 3
5 3 1 3 0 0
16 3 0 3 0 0 3 0 1 3 3 1 3 2 0 1 3
2 3 3
4 3 0 3 3
14 3 3 0 0 3 3 1 0 1 3 3 3 0 0
8 3 3 0 2 0 3 0 3
4 3 0 3 3
2 3 3
2 3 3
21 3 3 1 3 3 0 1 2 2 0 3 0 1 3 1 3 3 0 1 0 0
16 3 1 1 3 3 2 2 0 3 1 3 0 1 1 2 3
10 3 3 0 2 1 2 0 0 3 3
7 3 0 3 0 1 2 0
7 3 0 3 0 3 1 2
3 3 1 3
6 3 3 0 2 0 3
5 3 3 1 3 3
3 3 3 0
15 3 3 0 2 0 3 0 3 0 2 0 3 0 1 0
19 3 0 3 0 2 3 2 0 3 1 3 3 1 0 1 2 1 1 0
2 3 3
3 3 1 3
8 3 2 0 3 1 3 3 0
6 3 0 3 0 3 3
17 3 3 0 2 1 3 3 1 3 0 2 3 1 2 1 1 1
2 3 3
13 3 1 3 0 0 1 3 0 0 0 1 0 2
2 3 3
12 3 0 3 1 2 1 1 1 0 1 2 3
7 3 0 3 0 3 3 0
11 3 0 3 0 2 0 0 2 0 0 2
13 3 1 1 1 1 1 1 1 3 0 3 3 1
6 3 0 3 0 2 0
4 3 3 0 0
10 3 3 2 0 1 1 1 1 1 1
6 3 3 0 0 3 3
4 3 2 3 0
13 3 2 0 1 3 1 3 3 3 1 3 1 3
1 3
9 3 0 2 3 0 2 0 3 3
9 3 3 2 3 0 1 2 0 3
1 3
3 3 0 3
4 3 0 3 3
14 3 1 2 0 2 0 3 0 1 3 3 1 3 0
4 3 0 3 3
2 3 3
20 3 3 1 2 1 3 0 0 1 3 0 0 1 2 3 1 3 3 1 3
15 3 3 3 0 1 3 3 3 3 0 3 1 3 3 3
1 3
11 3 0 3 0 3 0 1 3 3 0 3
25 3 1 3 1 3 2 3 0 1 2 1 3 1 3 3 1 1 1 2 1 2 0 3 1 2
8 3 3 1 1 1 1 3 3
7 3 3 0 2 0 3 0
11 3 3 1 1 1 1 1 3 0 0 3
3 3 1 3
5 3 0 1 0 3
22 3 3 0 0 0 1 2 3 3 1 1 1 1 1 1 3 3 0 1 3 1 2
8 3 0 3 0 1 3 3 3
7 3 3 3 1 3 0 0
6 3 0 3 0 2 3
12 3 1 1 1 3 3 3 1 1 3 0 3
2 3 3
1 3
4 3 1 1 3
13 3 1 3 0 0 3 3 1 1 3 0 1 0
10 3 3 2 1 3 3 0 1 3 3
15 3 1 1 2 3 3 0 2 1 2 0 0 0 2 3
1 3
9 3 3 0 2 0 3 1 2 3
2 3 3
6 3 0 3 0 3 3
15 3 3 0 1 2 3 1 3 3 3 1 3 3 3 3
9 3 0 3 1 0 1 2 2 3
2 3 3
11 3 0 3 0 3 1 2 0 3 3 0
3 3 1 3
5 3 0 3 3 2
6 3 3 0 0 1 3
1 3
10 3 3 0 2 0 3 3 3 1 3
18 3 3 0 0 1 1 3 0 2 1 1 3 3 0 3 3 3 2
5 3 3 1 3 3
6 3 0 3 0 1 2
1 3
19 3 2 0 3 0 2 1 1 3 3 1 3 3 1 2 3 0 1 3
3 3 0 3
10 3 3 1 3 3 0 0 3 0 2
1 3
9 3 0 3 1 1 3 3 0 3
2 3 3
8 3 1 1 3 0 2 0 3
3 3 0 1
1 3
6 3 0 3 0 2 3
3 3 0 3
3 3 1 3
3 3 0 3
13 3 0 3 1 1 3 0 3 0 3 0 1 3
2 3 3
5 3 0 2 1 3
2 3 3
3 3 3 0
17 3 3 2 0 2 0 3 3 3 0 3 1 2 0 3 0 1
8 3 0 3 1 0 1 2 3
33 3 3 0 1 1 0 1 3 1 0 3 3 3 1 1 1 2 2 0 3 1 3 0 3 2 2 3 0 1 3 0 2 3
6 3 1 3 2 3 2
1 3
2 3 3
9 3 0 3 0 2 3 1 2 1
3 3 0 3
7 3 0 1 3 3 0 3
7 3 3 1 3 3 0 3
2 3 0
5 3 0 3 1 3
4 3 0 1 0
2 3 3
11 3 0 3 0 1 3 3 1 3 3 2
8 3 3 1 1 2 1 0 2
9 3 0 3 1 2 1 3 2 3
5 3 3 1 3 1
6 3 3 0 1 1 1
28 3 3 0 2 2 0 3 0 2 3 2 0 0 0 3 0 0 1 1 3 1 1 2 0 2 3 0 1
2 3 3
3 3 3 0
21 3 3 0 1 2 0 0 2 3 0 2 3 1 3 3 3 0 2 2 0 3
6 3 3 1 3 0 3
8 3 0 3 0 1 3 3 3
4 3 1 3 0
6 3 2 0 3 1 0
8 3 3 0 0 0 1 1 3
2 3 3
7 3 0 2 3 2 0 3
6 3 0 3 1 2 3
8 3 3 1 3 3 1 2 3
4 3 0 3 0
3 3 3 0
11 3 3 1 3 1 3 0 1 1 1 0
4 3 0 2 3
3 3 3 2
9 3 3 0 0 1 3 0 0 0
1 3
30 3 1 2 0 2 0 3 1 2 1 3 0 2 3 2 0 0 2 3 1 1 1 3 1 3 1 3 3 3 2
5 3 3 0 2 3
2 3 3
5 3 3 2 2 3
6 3 3 1 1 3 0
1 3
8 3 0 3 3 2 3 0 1
1 3
10 3 0 3 1 3 0 2 2 0 3
9 3 3 1 3 3 0 2 3 0
7 3 0 3 1 1 0 3
11 3 1 0 1 0 2 0 0 3 0 2
11 3 3 2 0 2 0 3 1 2 0 3
11 3 0 1 1 1 1 2 0 3 0 3
16 3 3 1 1 3 2 1 2 0 2 3 0 2 1 3 0
5 3 1 1 2 0
2 3 3
3 3 3 0
3 3 1 3
1 3
2 3 1
5 3 0 1 0 3
25 3 0 1 2 1 1 3 0 2 1 1 1 1 3 0 3 3 3 0 1 3 3 3 0 2
2 3 3
3 3 3 0
2 3 3
5 3 0 3 0 2
6 3 3 0 0 1 3
9 3 0 3 0 1 2 3 1 0
4 3 3 0 2
10 3 1 1 3 1 3 3 0 2 3
14 3 3 1 0 2 1 3 3 3 0 2 3 0 3
6 3 3 3 3 3 2
9 3 3 2 0 1 0 1 2 3
9 3 0 3 3 0 2 0 2 3
3 3 3 0
12 3 1 3 0 1 1 1 2 0 3 0 2
2 3 3
11 3 0 2 1 3 0 1 2 0 2 3
3 3 1 3
4 3 0 3 0
7 3 1 1 2 3 0 3
2 3 2
5 3 3 0 0 3
4 3 1 3 0
11 3 0 2 1 3 1 3 3 1 3 0
1 3
18 3 0 3 0 0 1 1 1 2 0 3 0 1 3 3 1 2 3
1 3
22 3 0 3 1 2 1 1 1 1 1 2 0 3 0 0 3 0 2 0 1 2 3
3 3 3 0
8 3 1 1 1 1 3 1 3
10 3 0 3 3 0 2 1 2 0 2
5 3 3 0 2 1
5 3 3 1 3 3
10 3 0 3 3 1 3 3 0 3 0
4 3 0 2 3
14 3 0 1 0 1 3 0 2 1 1 1 3 1 3
12 3 1 3 1 3 3 1 2 1 1 3 1
2 3 3
5 3 3 0 0 0
5 3 2 0 0 3
2 3 3
4 3 1 3 0
15 3 1 3 0 1 2 0 3 1 2 2 0 3 0 0
2 3 3
7 3 0 3 1 0 1 0
10 3 0 0 3 2 1 2 0 2 3
4 3 1 1 3
6 3 3 0 0 0 1
6 3 0 3 0 1 2
8 3 3 0 0 1 3 0 0
7 3 3 0 1 1 1 3
4 3 1 3 0
2 3 3
2 3 1
15 3 1 1 3 1 3 3 1 3 0 3 0 0 3 0
28 3 3 0 0 0 1 0 1 2 0 3 0 0 3 3 1 3 0 3 0 1 0 1 0 2 2 1 3
2 3 3
2 3 3
10 3 0 0 3 2 0 3 0 1 0
3 3 0 3
15 3 0 3 3 3 0 2 3 0 2 0 3 1 3 3
27 3 1 1 1 1 0 3 3 0 3 0 0 3 1 0 1 3 3 1 2 2 0 3 3 0 2 0
13 3 3 3 1 3 3 0 3 0 1 0 0 2
10 3 3 1 3 3 0 3 1 2 3
21 3 0 3 0 2 3 1 2 2 0 3 0 0 3 0 1 3 3 1 3 0
5 3 0 2 1 3
2 3 3
7 3 1 3 1 3 0 2
14 3 3 1 3 3 0 3 0 0 1 3 3 0 3
12 3 1 1 1 1 1 1 3 0 3 3 3
17 3 3 1 3 3 0 1 3 3 0 3 0 3 0 1 2 1
1 3
3 3 0 3
23 3 0 3 1 2 3 1 3 3 1 3 3 0 3 3 1 0 1 2 2 0 3 0
2 3 0
3 3 0 3
2 3 3
4 3 1 3 0
2 3 3
6 3 3 1 3 0 0
3 3 0 3
4 3 3 2 3
4 3 0 2 3
3 3 3 1
7 3 3 0 0 1 3 0
1 3
2 3 3
4 3 0 3 3
1 3
11 3 0 3 1 0 2 0 1 3 0 3
3 3 1 0
11 3 3 0 1 1 1 0 3 2 2 3
8 3 0 3 1 0 1 3 3
3 3 0 3
3 3 3 0
10 3 3 0 0 3 3 3 3 3 0
4 3 3 2 0
4 3 1 1 3
8 3 0 3 1 2 2 0 3
1 3
3 3 3 0
5 3 3 0 2 1
15 3 0 3 0 3 0 2 0 3 1 1 1 1 3 0
14 3 3 0 0 1 3 0 0 1 3 0 2 0 1
1 3
1 3
3 3 0 3
8 3 3 2 0 0 1 0 2
7 3 0 2 1 3 0 0
13 3 3 0 2 0 3 0 1 0 1 3 3 3
2 3 3
8 3 3 2 1 0 1 3 3
2 3 3
2 3 3
6 3 3 1 3 3 3
7 3 1 3 1 3 3 3
1 3
1 3
25 3 0 3 3 1 3 3 0 3 0 0 3 0 1 0 2 2 2 3 0 2 1 3 2 1
1 3
9 3 3 1 3 3 0 1 0 3
2 3 3
1 3
9 3 0 3 3 0 0 1 1 3
6 3 1 3 0 0 3
15 3 0 3 3 1 3 3 1 1 3 0 1 0 0 0
7 3 0 3 3 1 0 0
4 3 3 0 2
3 3 1 3
1 3
8 3 1 3 1 0 3 3 0
4 3 0 2 3
8 3 3 1 3 3 1 3 0
8 3 3 3 1 3 3 0 2
6 3 3 0 1 0 2
3 3 1 1
7 3 0 3 2 0 1 3
9 3 3 3 0 2 3 1 3 0
3 3 0 3
3 3 3 0
21 3 0 3 0 2 2 2 3 0 2 0 3 1 3 3 1 3 3 3 2 0
11 3 3 3 3 1 3 0 0 2 0 3
2 3 3
7 3 1 1 3 3 3 2
4 3 0 3 3
14 3 2 0 3 0 2 0 3 0 2 0 1 3 0
7 3 3 1 3 3 0 3
1 3
6 3 0 3 1 3 0
10 3 0 2 3 3 0 3 3 3 0
4 3 0 2 0
4 3 1 3 2
7 3 2 0 3 1 3 3
3 3 0 3
10 3 3 1 3 3 0 1 3 3 3
4 3 1 3 0
1 3
2 3 3
3 3 0 3
2 3 3
7 3 0 1 2 2 0 1
19 3 2 0 3 1 3 2 3 0 2 3 0 1 2 3 0 0 1 3
4 3 3 1 2
3 3 3 0
7 3 3 0 0 1 3 0
5 3 0 0 2 3
4 3 1 1 2
2 3 3
5 3 0 3 0 2
6 3 3 0 1 2 3
3 3 0 3
3 3 0 2
1 3
7 3 3 1 3 3 1 3
13 3 0 3 3 0 1 2 3 0 2 0 3 0
1 3
5 3 0 2 3 0
7 3 1 3 1 3 0 3
3 3 3 2
6 3 1 3 1 1 1
7 3 0 3 0 1 3 3
3 3 0 3
1 3
19 3 0 3 1 0 1 3 3 0 3 0 1 3 0 0 0 1 3 3
1 3
9 3 0 0 0 1 3 3 3 0
5 3 0 3 1 2
3 3 3 2
7 3 3 1 3 3 0 3
5 3 3 0 0 0
3 3 1 3
4 3 0 2 3
2 3 3
6 3 0 3 1 3 0
5 3 0 1 0 0
3 3 0 3
6 3 3 0 2 3 3
8 3 3 2 0 1 3 1 2
6 3 3 0 0 1 3
3 3 3 3
4 3 2 0 3
3 3 0 3
4 3 1 1 3
14 3 3 1 3 3 3 1 3 3 0 3 0 1 0
7 3 1 3 0 0 0 3
2 3 3
7 3 3 1 3 1 0 3
3 3 1 3
23 3 3 1 3 3 1 2 1 2 0 3 0 0 1 1 1 2 0 3 1 2 3 0
6 3 3 1 2 3 3
5 3 3 0 1 3
4 3 1 1 3
6 3 1 2 0 1 3
4 3 1 1 2
7 3 0 3 1 3 0 3
1 3
2 3 3
5 3 0 2 1 3
3 3 1 3
7 3 0 3 1 2 1 3
10 3 0 1 2 0 3 3 0 2 2
14 3 3 0 3 3 0 3 0 3 0 2 0 0 2
7 3 1 3 3 3 0 2
5 3 0 3 0 2
4 3 3 1 1
4 3 3 0 2
14 3 0 3 1 0 1 2 3 1 1 3 0 3 3
9 3 0 3 1 0 1 3 3 3
3 3 0 3
4 3 2 0 3
9 3 1 1 3 3 0 1 3 3
2 3 3
7 3 0 3 1 2 3 3
2 3 3
6 3 3 0 2 0 3
3 3 3 1
7 3 3 1 3 3 3 2
4 3 1 3 0
9 3 0 3 0 3 1 3 1 3
4 3 1 3 0
4 3 2 0 3
4 3 1 3 0
2 3 3
9 3 0 3 1 0 1 3 3 3
24 3 0 3 1 3 2 0 3 0 0 3 3 1 1 1 1 1 1 3 3 2 0 0 3
13 3 0 3 0 1 3 3 1 3 0 2 0 3
3 3 0 3
5 3 0 3 3 0
1 3
4 3 0 3 3
2 3 3
6 3 1 0 3 3 0
2 3 0
7 3 3 3 1 3 3 0
13 3 3 3 1 2 3 3 1 2 3 1 3 3
5 3 3 1 3 3
28 3 0 3 1 2 2 0 3 1 2 2 2 1 1 1 1 3 3 1 0 0 2 3 1 1 1 3 0
5 3 1 1 1 3
4 3 0 3 0
2 3 3
8 3 3 1 3 3 1 3 3
7 3 3 1 0 1 0 0
15 3 0 3 0 0 1 2 1 2 1 1 3 3 3 0
14 3 3 0 1 2 3 1 3 3 1 2 0 3 0
3 3 0 3
4 3 1 2 2
19 3 2 0 1 1 3 0 2 3 1 3 3 1 1 1 1 2 3 1
1 3
4 3 1 3 0
17 3 0 3 0 1 2 3 0 2 3 1 3 2 2 3 0 3
9 3 0 1 3 3 1 0 0 0
4 3 0 3 3
2 3 3
25 3 1 1 3 0 0 3 0 1 3 3 0 1 2 3 0 0 3 3 1 0 1 2 1 0
5 3 0 3 1 3
16 3 0 3 0 3 0 0 3 1 3 3 0 2 2 0 3
2 3 3
7 3 1 3 1 3 0 2
1 3
7 3 3 1 3 0 1 0
6 3 3 0 0 1 3
3 3 1 3
27 3 2 0 3 1 3 2 0 1 3 3 3 0 2 3 3 1 3 0 2 2 0 3 0 2 0 3
11 3 1 3 0 2 1 1 3 3 3 0
3 3 1 3
8 3 3 1 3 3 3 2 0
8 3 1 1 3 0 0 1 3
4 3 0 3 3
9 3 3 0 2 1 0 3 3 3
22 3 1 1 3 0 1 1 2 0 3 0 1 3 3 0 1 3 3 1 0 1 3
9 3 3 0 1 1 1 3 2 2
9 3 3 1 3 3 1 3 3 2
11 3 0 1 3 3 0 1 2 3 3 0
11 3 3 1 2 3 0 3 0 2 3 1
21 3 1 3 0 1 0 2 3 2 0 1 2 2 3 1 3 3 1 3 0 3
27 3 3 1 3 2 0 1 3 3 0 1 3 3 0 3 0 2 1 1 3 3 0 1 1 2 0 3
5 3 0 3 1 3
2 3 0
4 3 3 0 0
1 3
3 3 0 3
6 3 3 0 2 1 3
8 3 3 0 2 1 1 2 0
3 3 0 3
11 3 3 0 2 0 3 0 1 3 3 3
3 3 3 0
3 3 1 3
2 3 0
3 3 1 3
7 3 1 3 0 0 1 3
3 3 0 3
4 3 0 3 0
4 3 0 3 3
6 3 0 3 1 3 1
8 3 0 2 3 0 0 1 3
22 3 0 2 3 1 3 3 1 3 0 3 1 2 1 1 2 3 1 3 3 1 2
3 3 0 2
8 3 0 3 1 0 1 3 2
2 3 3
3 3 0 3
10 3 0 0 1 3 0 3 0 3 3
9 3 0 3 0 3 3 3 3 0
31 3 2 0 3 0 2 1 2 0 2 0 3 0 1 3 3 1 2 0 3 0 2 0 3 0 1 3 3 1 3 0
1 3
5 3 0 3 3 3
4 3 0 1 1
4 3 3 0 3
3 3 0 3
3 3 3 2
4 3 0 3 0
11 3 0 3 0 1 1 3 1 1 3 0
14 3 0 3 1 2 0 1 3 0 2 1 0 3 3
19 3 0 3 0 3 3 2 2 3 3 3 3 1 3 3 1 2 1 3
3 3 0 3
1 3
5 3 1 0 3 2
5 3 3 0 0 0
1 3
2 3 3
7 3 0 3 0 1 3 3
2 3 3
7 3 0 2 3 0 0 0
1 3
19 3 1 0 3 0 2 3 1 1 3 0 3 2 1 1 0 1 0 0
2 3 1
17 3 1 1 3 3 1 1 3 0 1 2 3 0 0 1 3 0
10 3 0 3 1 0 2 3 0 2 3
4 3 1 1 3
5 3 1 3 3 0
3 3 0 3
3 3 0 3
2 3 3
1 3
4 3 0 1 0
6 3 2 0 0 3 0
5 3 0 2 3 0
10 3 0 3 0 3 3 0 2 0 3
4 3 1 3 1
4 3 1 3 0
6 3 3 0 0 1 3
1 3
21 3 2 0 0 3 0 1 1 2 0 3 1 2 0 3 0 0 3 3 0 3
1 3
12 3 3 1 3 3 3 0 0 3 3 0 3
25 3 0 3 0 1 2 3 1 3 0 2 1 3 1 3 2 2 0 3 0 2 3 2 0 3
12 3 1 3 0 0 0 1 1 0 2 3 2
2 3 3
1 3
4 3 1 3 0
4 3 0 3 3
22 3 0 3 1 2 2 1 3 0 2 1 1 0 3 3 1 0 3 3 3 2 3
5 3 1 0 3 0
17 3 0 3 1 2 1 3 1 3 3 3 3 0 2 0 2 3
10 3 0 3 0 1 1 1 3 1 3
5 3 2 0 3 1
3 3 3 0
1 3
6 3 3 0 2 0 3
4 3 3 0 2
2 3 3
27 3 0 3 1 2 1 1 3 2 2 3 2 3 1 1 3 0 3 0 1 3 3 1 3 1 1 2
2 3 2
1 3
1 3
5 3 0 1 2 3
2 3 3
3 3 0 3
3 3 0 3
2 3 3
18 3 0 3 0 1 0 1 3 3 3 1 3 3 1 3 0 2 3
1 3
4 3 1 3 3
4 3 0 3 2
3 3 0 3
9 3 0 1 3 3 1 1 3 0
2 3 0
8 3 3 0 2 0 3 0 2
4 3 0 2 3
4 3 0 3 1
2 3 3
15 3 1 1 1 1 1 2 0 3 1 2 1 1 1 1
4 3 3 0 0
3 3 3 1
6 3 0 3 0 3 0
10 3 3 1 3 3 1 3 3 0 1
4 3 0 3 3
2 3 1
7 3 0 2 3 3 1 3
6 3 1 3 1 1 1
4 3 0 2 3
3 3 3 0
4 3 1 1 3
5 3 0 2 1 3
3 3 3 2
2 3 0
7 3 3 0 2 2 0 3
8 3 3 1 3 3 0 3 3
2 3 3
9 3 3 0 2 1 3 3 0 0
6 3 0 3 1 3 3
27 3 0 3 1 1 3 3 3 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0
3 3 0 1
4 3 1 3 0
2 3 3
7 3 1 1 3 1 2 0
7 3 3 1 3 3 0 1
10 3 3 3 0 2 2 0 3 1 0
7 3 3 2 0 1 3 2
9 3 0 3 1 0 1 3 3 2
3 3 3 2
2 3 0
5 3 0 3 3 0
11 3 0 3 1 3 3 1 1 3 3 2
5 3 3 0 0 0
6 3 3 0 1 1 1
6 3 3 3 1 3 1
2 3 0
2 3 3
5 3 0 2 3 0
10 3 3 0 2 0 3 1 3 3 2
4 3 1 3 0
9 3 3 1 3 3 1 2 1 0
4 3 2 0 3
3 3 0 3
7 3 0 3 0 1 3 3
3 3 1 2
3 3 0 3
6 3 0 3 0 1 1
3 3 3 2
1 3
4 3 1 1 1
1 3
2 3 3
3 3 1 3
2 3 3
15 3 3 1 3 3 3 2 2 3 0 2 0 1 1 3
7 3 3 1 2 0 0 2
6 3 0 3 3 1 1
6 3 3 0 1 2 3
3 3 0 3
5 3 1 3 3 2
6 3 0 3 1 2 3
3 3 1 3
6 3 3 1 1 1 3
2 3 3
3 3 3 0
4 3 0 1 2
2 3 3
4 3 0 2 3
5 3 1 3 0 1
1 3
5 3 0 2 1 3
3 3 1 2
19 3 3 1 3 3 2 1 1 1 0 1 3 3 3 1 1 3 0 0
10 3 0 3 0 0 3 2 0 3 0
14 3 0 3 0 1 3 3 1 3 0 2 0 3 0
2 3 3
4 3 0 3 2
17 3 0 3 0 1 3 3 1 2 1 2 1 1 3 3 1 3
12 3 3 3 0 1 1 1 1 1 1 1 1
3 3 1 3
20 3 0 1 1 2 3 0 2 1 1 3 3 3 1 0 1 3 3 0 3
29 3 1 3 0 1 1 2 0 3 1 3 1 1 1 2 3 0 1 3 1 1 1 2 1 0 0 0 1 2
6 3 1 1 3 0 2
3 3 3 1
5 3 3 0 1 3
11 3 0 3 1 2 3 0 2 2 0 3
10 3 3 0 2 0 3 1 2 1 1
57 3 0 3 0 3 0 2 0 0 0 1 1 3 3 1 1 3 0 1 1 1 1 1 1 1 1 2 3 1 3 3 1 2 1 0 1 2 0 2 3 0 3 1 3 0 2 1 0 2 0 0 0 1 3 0 0 0
2 3 3
7 3 1 3 0 1 1 3
3 3 0 3
11 3 0 3 0 3 0 1 3 3 0 2
5 3 1 3 3 3
13 3 3 0 1 3 2 2 0 3 1 1 3 3
12 3 1 1 3 3 0 3 0 1 3 3 3
5 3 1 1 3 0
14 3 1 2 1 3 3 0 3 0 1 3 3 3 0
2 3 3
13 3 0 1 1 3 1 3 0 2 3 3 0 0
3 3 3 1
3 3 0 3
4 3 0 2 3
3 3 3 0
2 3 3
1 3
9 3 3 1 1 1 2 0 3 3
9 3 0 2 3 0 1 2 1 3
6 3 3 1 3 3 3
26 3 3 0 1 2 0 3 0 3 0 1 3 3 3 1 2 3 1 3 1 3 3 0 2 0 3
2 3 3
7 3 0 3 0 0 3 0
3 3 0 2
2 3 1
2 3 3
5 3 3 1 0 2
8 3 3 0 2 3 2 0 2
6 3 0 3 0 3 0
5 3 0 2 3 0
9 3 3 1 2 2 1 3 0 1
1 3
6 3 0 1 0 2 0
11 3 0 1 3 3 3 3 0 2 1 2
5 3 1 3 0 0
9 3 3 1 3 3 0 2 3 0
6 3 0 3 3 2 3
3 3 1 1
4 3 2 0 3
5 3 0 2 3 1
4 3 0 3 3
2 3 0
4 3 3 2 0
2 3 3
13 3 3 2 0 2 0 3 1 3 2 0 3 0
5 3 0 3 0 2
5 3 0 3 1 0
9 3 0 3 0 3 3 1 3 3
33 3 3 2 2 2 3 0 0 0 3 3 3 0 1 3 3 0 2 0 0 2 1 3 2 0 2 0 3 1 3 0 3 3
5 3 3 1 3 3
11 3 3 3 2 3 0 2 2 0 3 0
10 3 0 3 0 2 3 3 3 0 2
11 3 0 3 0 1 3 3 0 3 3 0
6 3 0 3 1 2 3
4 3 3 1 2
4 3 1 1 3
9 3 1 3 0 1 3 2 0 3
19 3 3 0 1 1 1 1 3 3 3 3 0 2 1 3 0 0 1 3
2 3 1
3 3 0 3
2 3 3
4 3 0 3 3
4 3 2 0 3
11 3 0 3 0 3 1 1 1 1 3 0
5 3 1 3 0 2
4 3 1 2 3
5 3 2 0 3 0
8 3 0 3 0 0 1 3 3
8 3 1 0 3 3 0 1 2
3 3 1 3
5 3 3 0 2 3
5 3 0 3 3 0
5 3 0 3 3 2
4 3 3 2 3
10 3 0 3 1 0 1 3 3 1 0
4 3 0 3 0
7 3 3 1 2 2 1 3
5 3 0 3 3 0
6 3 0 3 2 0 3
6 3 0 2 1 1 3
3 3 0 3
3 3 1 2
6 3 3 0 2 1 0
8 3 0 3 0 1 3 2 0
9 3 1 3 0 2 2 0 3 0
20 3 2 3 0 1 3 3 0 1 1 3 3 3 0 3 0 2 2 0 3
7 3 3 3 0 0 0 2
17 3 3 0 1 0 1 3 3 3 0 1 3 3 0 3 1 3
13 3 0 3 3 1 3 3 0 1 2 3 0 2
5 3 1 3 0 2
9 3 0 3 3 2 3 3 3 3
10 3 0 3 2 0 3 0 1 3 1
20 3 1 3 1 3 0 2 0 3 1 3 0 2 0 3 0 2 3 0 2
3 3 0 3
2 3 0
8 3 0 3 0 3 0 3 3
3 3 0 3
9 3 0 3 0 2 0 0 1 2
17 3 3 0 0 3 3 1 2 2 0 3 0 3 1 2 0 3
19 3 1 3 1 3 0 2 3 3 2 3 1 3 0 3 0 3 0 2
12 3 3 1 0 2 1 1 2 2 0 3 0
10 3 3 0 0 1 3 1 3 1 0
4 3 1 2 0
4 3 1 3 0
20 3 0 3 0 1 3 3 0 3 0 1 3 3 3 0 1 1 2 0 3
4 3 0 1 1
6 3 0 3 3 1 0
2 3 3
8 3 0 3 1 2 2 0 1
4 3 1 3 0
10 3 3 0 1 0 1 3 3 0 0
1 3
4 3 3 0 0
4 3 3 1 2
12 3 3 1 3 3 0 3 3 1 3 2 3
2 3 0
7 3 3 1 3 3 3 1
4 3 1 3 0
1 3
3 3 0 3
3 3 3 2
2 3 3
4 3 1 0 3
1 3
33 3 1 3 2 0 2 0 2 0 0 1 3 3 0 1 3 0 1 3 3 3 3 0 2 0 3 0 3 1 3 3 0 0
23 3 1 3 0 0 3 3 1 3 0 3 0 2 3 3 1 3 0 1 1 1 0 1
4 3 1 0 0
3 3 0 3
8 3 0 3 1 2 1 1 3
5 3 1 3 0 0
8 3 3 2 1 3 3 1 3
16 3 1 3 1 3 3 0 3 1 2 1 1 0 1 3 2
4 3 1 3 0
13 3 0 3 0 1 3 3 0 2 2 1 1 1
6 3 0 3 0 1 0
5 3 3 0 0 0
3 3 0 2
20 3 0 3 0 2 0 1 0 1 2 1 0 0 2 3 0 2 0 3 0
4 3 1 1 3
4 3 3 0 2
3 3 0 3
8 3 2 3 0 2 0 1 3
15 3 1 3 0 3 3 3 0 2 0 2 3 0 1 0
4 3 0 3 3
21 3 3 0 1 1 1 2 0 3 1 0 1 3 3 0 3 1 3 0 3 0
7 3 0 3 1 2 1 0
6 3 0 3 0 2 3
14 3 0 3 0 1 3 3 0 3 3 0 2 0 2
1 3
2 3 3
10 3 0 3 0 0 3 1 0 2 0
29 3 3 1 3 3 0 3 0 3 3 1 0 2 1 1 1 2 0 2 0 0 2 1 2 0 1 2 3 0
3 3 3 0
8 3 0 2 3 0 0 1 3
20 3 0 3 1 2 1 3 1 0 1 3 3 1 0 1 3 3 1 3 0
6 3 1 3 0 2 3
15 3 0 3 3 0 0 1 3 1 0 3 3 0 3 0
2 3 3
5 3 1 1 3 3
26 3 1 3 1 1 1 1 1 1 1 1 3 3 3 0 2 1 1 3 0 0 1 1 3 0 2
3 3 3 2
10 3 0 3 1 2 1 1 3 0 2
5 3 3 0 1 1
4 3 0 2 3
5 3 0 3 0 2
12 3 0 3 3 2 3 1 1 3 0 3 0
2 3 3
2 3 3
4 3 3 0 2
5 3 3 3 1 3
15 3 0 3 1 2 1 2 1 3 3 0 3 3 3 3
9 3 3 0 2 1 1 3 0 1
6 3 0 3 0 3 3
2 3 3
11 3 0 3 1 3 0 3 1 3 0 1
9 3 1 3 0 0 1 1 1 3
2 3 3
11 3 1 2 0 0 1 1 3 0 1 0
5 3 3 0 1 3
2 3 3
5 3 3 1 3 3
4 3 3 0 1
4 3 0 3 3
6 3 1 1 3 1 3
1 3
12 3 3 3 1 3 3 3 0 0 1 3 0
16 3 1 1 3 0 0 0 3 0 0 2 3 2 2 0 2
4 3 3 0 0
9 3 0 3 1 2 2 0 3 3
6 3 0 3 0 2 3
6 3 3 1 3 0 2
7 3 0 3 1 2 0 3
3 3 1 2
7 3 1 3 0 1 1 0
6 3 0 2 3 0 0
5 3 3 1 1 3
9 3 0 3 1 3 1 3 3 3
15 3 2 0 3 0 2 0 3 0 0 1 3 3 1 3
10 3 3 0 1 1 2 3 3 2 0
4 3 1 1 3
3 3 1 3
9 3 0 3 3 1 3 3 0 2
6 3 3 2 0 0 2
2 3 0
10 3 0 2 0 0 0 1 3 0 0
5 3 0 3 1 3
1 3
67 3 3 3 0 1 3 2 1 3 2 0 2 3 2 0 3 1 0 1 2 1 1 1 1 2 0 3 0 3 1 3 0 3 1 2 0 3 3 1 3 3 3 0 1 3 2 3 0 2 2 0 3 0 1 1 2 3 1 2 0 1 3 0 0 1 3 0
4 3 0 3 0
3 3 0 3
4 3 1 3 0
3 3 3 2
2 3 3
16 3 0 3 0 3 0 1 3 3 3 3 0 0 3 0 0
2 3 3
2 3 3
4 3 3 0 0
15 3 1 3 3 1 3 1 2 3 1 1 0 2 0 3
6 3 0 2 1 1 3
7 3 0 1 3 3 3 0
3 3 0 3
8 3 0 3 1 3 3 0 0
2 3 3
16 3 1 1 3 1 1 3 1 1 1 1 3 3 3 0 3
3 3 1 1
2 3 3
18 3 3 2 3 0 3 0 2 3 0 3 1 2 1 1 0 0 3
19 3 3 1 3 0 2 3 1 3 1 3 3 1 0 1 0 1 0 0
3 3 0 3
3 3 1 3
28 3 0 3 1 2 0 1 0 1 3 0 2 2 3 1 3 3 0 1 3 3 0 0 2 0 3 1 3
3 3 0 3
3 3 0 3
2 3 3
4 3 0 1 0
3 3 1 3
4 3 3 3 2
3 3 1 3
15 3 1 3 0 2 1 1 3 0 0 2 1 3 0 1
2 3 3
20 3 0 2 3 0 1 3 2 0 3 0 0 1 3 1 3 3 1 2 3
6 3 3 1 3 0 3
3 3 1 3
18 3 1 2 0 0 3 3 0 3 0 2 1 2 0 0 1 3 0
2 3 3
2 3 3
2 3 0
8 3 0 3 3 0 2 0 3
17 3 1 3 0 2 2 2 3 3 3 3 3 3 2 3 0 3
28 3 0 0 2 3 0 1 1 2 0 3 0 1 3 3 1 0 1 3 3 1 2 0 3 0 1 2 3
7 3 3 1 3 3 0 3
1 3
2 3 3
10 3 3 1 3 3 3 1 2 3 3
1 3
3 3 3 0
20 3 3 1 3 3 0 2 0 3 0 2 1 3 2 0 2 1 1 1 1
15 3 0 3 1 2 2 0 3 0 1 1 3 3 3 2
10 3 0 2 3 0 2 0 1 0 0
17 3 0 3 1 0 2 0 2 1 1 3 3 3 3 1 2 3
11 3 3 1 0 3 0 0 1 2 1 3
4 3 1 1 3
2 3 3
9 3 0 3 1 2 1 1 2 0
6 3 1 3 0 2 3
10 3 3 0 1 0 3 0 1 1 3
12 3 3 0 2 3 1 3 3 3 3 0 2
5 3 0 3 3 0
6 3 0 3 2 0 3
16 3 0 3 1 2 1 0 2 2 0 1 3 0 2 3 0
6 3 3 0 2 1 2
7 3 3 3 1 3 0 0
9 3 1 1 1 3 1 3 3 3
9 3 0 3 1 0 3 3 3 0
6 3 1 1 3 0 0
7 3 3 1 3 3 1 0
3 3 3 2
3 3 0 3
4 3 0 2 3
6 3 0 0 2 0 3
11 3 0 1 3 3 1 3 0 0 0 1
9 3 3 0 0 0 3 3 3 3
8 3 3 1 0 0 1 0 0
3 3 3 0
7 3 0 3 0 0 2 3
8 3 0 2 3 0 2 1 2
5 3 0 2 3 3
2 3 3
1 3
13 3 3 1 3 0 0 2 0 3 0 1 2 1
4 3 3 0 2
2 3 3
9 3 0 2 3 1 0 1 1 3
12 3 3 1 2 2 0 3 1 2 0 3 0
3 3 3 0
14 3 1 3 1 1 1 3 0 0 0 3 3 3 3
26 3 1 0 2 3 0 2 0 3 0 1 3 3 0 2 3 0 1 2 3 2 1 0 1 3 3
5 3 0 3 0 3
4 3 2 0 3
10 3 3 3 2 0 0 1 3 3 3
23 3 0 1 2 1 2 3 0 0 1 3 0 1 2 0 3 0 1 3 3 0 1 0
7 3 1 3 0 1 1 3
8 3 0 2 3 1 3 3 3
12 3 0 3 0 3 1 3 1 1 3 0 0
15 3 3 0 0 0 3 3 3 0 1 3 3 0 0 3
10 3 3 3 0 1 1 1 1 1 3
9 3 0 3 3 0 2 2 0 3
7 3 0 3 0 3 1 2
3 3 3 0
1 3
1 3
7 3 0 3 0 1 2 1
2 3 3
9 3 0 2 3 0 0 1 3 0
3 3 3 0
16 3 1 1 1 1 1 3 0 1 3 0 3 1 0 3 3
10 3 3 0 2 3 1 2 3 1 3
3 3 0 3
8 3 3 1 3 3 0 2 3
5 3 3 0 2 1
7 3 0 2 3 1 3 1
9 3 0 2 3 0 1 2 0 3
3 3 1 2
3 3 0 3
2 3 3
3 3 3 2
10 3 3 3 0 2 2 0 0 3 0
14 3 0 3 1 2 1 1 1 2 3 0 1 0 0
8 3 0 3 0 3 3 2 0
8 3 3 0 2 3 1 3 3
8 3 0 3 1 1 1 3 0
2 3 0
4 3 1 3 0
4 3 1 3 1
4 3 3 2 1
24 3 0 3 0 3 0 2 0 1 3 0 2 1 3 3 2 2 3 1 1 3 2 1 3
3 3 1 3
1 3
10 3 0 3 3 2 2 2 3 0 0
7 3 0 3 3 1 2 1
3 3 2 1
4 3 1 3 0
3 3 3 0
2 3 3
3 3 3 2
5 3 1 1 3 1
19 3 0 3 0 3 0 1 3 3 0 1 3 3 0 3 0 2 3 0
4 3 3 0 2
15 3 3 1 3 3 0 1 0 3 3 3 3 2 0 3
2 3 3
8 3 3 1 3 3 3 3 0
5 3 0 2 3 0
2 3 3
2 3 3
10 3 1 2 1 3 0 3 3 3 0
5 3 0 3 3 0
11 3 0 2 3 1 1 1 3 1 3 0
3 3 3 0
2 3 3
2 3 3
21 3 0 3 1 2 1 1 2 0 3 1 2 3 0 1 3 0 1 3 3 0
14 3 1 3 1 3 3 0 1 1 1 2 0 3 3
4 3 1 1 2
2 3 2
5 3 1 1 3 0
5 3 1 3 0 2
7 3 3 0 2 0 3 0
5 3 0 3 0 2
4 3 1 3 1
9 3 0 3 3 1 2 3 3 0
7 3 0 3 0 2 0 3
1 3
2 3 3
16 3 0 3 0 1 2 2 3 1 3 3 3 0 2 3 3
2 3 3
1 3
4 3 0 3 3
3 3 3 3
3 3 3 1
4 3 1 1 3
18 3 3 3 0 3 3 3 2 3 0 1 3 3 3 1 2 1 3
13 3 0 3 0 1 1 1 1 0 3 3 0 3
8 3 0 3 1 3 1 3 1
10 3 0 1 3 3 0 3 0 3 0
20 3 2 0 3 0 0 0 2 0 3 1 0 1 3 3 0 3 0 2 3
13 3 0 3 0 3 1 3 1 0 1 3 0 3
2 3 3
18 3 3 0 1 0 1 2 1 1 3 1 0 1 0 1 3 2 0
10 3 3 0 0 1 3 0 0 1 3
4 3 2 0 3
10 3 1 1 3 3 1 1 3 0 2
7 3 3 0 1 2 1 3
8 3 1 1 3 3 0 1 0
19 3 0 3 3 0 2 0 3 1 3 3 0 1 0 1 3 3 0 2
7 3 0 3 1 3 0 3
9 3 3 1 3 3 2 1 3 3
50 3 2 0 3 0 2 1 1 3 3 0 3 0 3 3 0 2 1 2 0 0 1 3 1 3 3 1 2 0 1 3 3 0 2 0 3 1 0 1 3 3 1 0 3 3 0 3 1 2 1
4 3 1 3 0
13 3 0 3 0 1 0 0 1 1 0 1 3 0
4 3 3 2 2
2 3 3
2 3 3
7 3 3 0 2 0 3 0
20 3 3 3 1 3 3 1 2 0 3 0 0 3 3 3 3 3 0 0 3
7 3 3 1 3 3 1 3
9 3 3 1 3 3 2 0 1 3
4 3 0 0 3
12 3 0 3 3 1 0 1 3 3 2 0 3
10 3 3 0 1 2 0 3 1 3 3
8 3 0 3 0 3 1 1 3
7 3 0 3 1 3 3 0
7 3 3 1 3 3 0 3
5 3 2 0 1 3
14 3 0 3 1 2 1 2 3 1 3 3 1 0 2
9 3 3 1 1 1 2 0 2 3
16 3 0 0 2 1 1 0 0 3 0 2 0 1 1 3 0
2 3 3
10 3 0 3 1 2 1 1 2 0 3
14 3 0 3 3 1 3 3 0 3 1 1 3 0 1
4 3 1 1 3
18 3 0 3 1 3 0 0 1 3 0 0 1 3 0 2 0 3 0
9 3 3 2 1 3 3 1 3 3
16 3 3 1 1 3 0 1 3 3 1 2 3 0 2 0 3
3 3 0 3
12 3 0 3 3 1 2 1 1 1 1 1 3
3 3 1 3
6 3 0 2 3 0 2
7 3 0 3 0 1 3 3
10 3 3 1 3 3 1 3 2 0 3
13 3 1 1 1 1 3 0 2 0 1 2 3 0
5 3 3 1 3 3
2 3 3
3 3 1 3
11 3 1 1 3 3 3 1 1 0 2 1
6 3 0 3 1 3 3
9 3 0 3 0 3 0 1 3 1
4 3 0 1 0
17 3 3 0 0 1 3 0 0 0 2 1 3 1 3 1 3 3
4 3 1 3 0
3 3 3 0
26 3 3 2 1 3 3 0 3 0 1 3 3 0 3 1 3 0 3 1 3 3 1 1 3 2 3
8 3 3 0 0 0 3 3 3
6 3 3 0 0 3 3
13 3 0 3 3 0 1 2 1 3 0 1 2 3
6 3 3 2 0 1 3
1 3
17 3 1 3 1 1 1 3 3 2 1 1 2 0 3 0 3 3
2 3 3
6 3 3 0 1 1 1
21 3 0 3 0 1 2 0 3 0 2 1 2 0 0 1 3 0 2 0 3 0
13 3 0 3 1 2 1 2 3 1 3 1 3 0
10 3 0 3 0 2 3 1 1 3 3
3 3 0 3
10 3 0 3 1 3 0 2 2 0 3
3 3 0 3
3 3 3 2
4 3 0 3 0
26 3 3 1 3 3 0 1 3 3 0 1 3 3 1 2 2 3 1 3 3 3 0 1 2 1 3
6 3 0 3 3 0 2
7 3 3 0 0 0 1 0
9 3 0 2 1 3 0 2 1 0
5 3 0 3 1 3
9 3 3 2 0 2 1 3 0 1
2 3 0
27 3 1 1 3 3 3 0 2 0 3 1 2 3 0 2 1 0 3 3 3 1 3 3 3 0 2 0
8 3 3 0 3 3 0 3 1
5 3 1 3 0 2
12 3 0 3 0 3 3 0 1 3 2 1 0
21 3 0 1 2 1 1 3 0 3 1 3 3 1 3 3 1 3 3 3 0 3
1 3
3 3 0 3
6 3 0 3 1 2 3
4 3 3 1 3
3 3 1 3
3 3 3 0
24 3 1 1 3 0 1 1 1 1 3 1 3 3 3 0 2 3 0 3 0 1 3 3 3
13 3 2 0 3 1 1 3 2 3 0 0 3 3
9 3 2 0 1 3 0 2 0 3
6 3 0 1 0 3 2
2 3 3
3 3 0 3
12 3 0 3 0 3 1 3 3 3 1 3 0
14 3 3 2 0 1 3 0 3 0 3 0 3 3 3
3 3 3 0
5 3 0 3 0 1
1 3
4 3 1 2 0
5 3 3 1 3 3
8 3 3 0 1 0 3 0 2
3 3 0 1
7 3 0 3 2 0 1 3
7 3 3 0 2 0 1 0
3 3 3 1
1 3
7 3 0 3 1 3 3 3
6 3 3 3 1 3 3
3 3 0 3
16 3 0 3 1 1 3 3 0 1 2 0 1 3 3 1 3
2 3 3
14 3 3 1 0 0 2 1 2 0 3 0 3 1 2
3 3 0 3
10 3 1 1 3 1 3 0 2 0 2
2 3 0
14 3 1 2 0 0 3 3 1 3 3 1 1 1 1
9 3 0 2 3 0 1 2 3 2
15 3 0 3 0 0 1 2 3 0 1 2 1 2 1 3
13 3 3 1 3 3 1 3 3 3 3 0 1 3
10 3 3 0 2 1 1 1 1 2 0
1 3
6 3 0 3 1 3 3
3 3 0 3
3 3 0 1
2 3 0
6 3 3 2 1 2 2
6 3 3 1 3 3 0
3 3 0 3
7 3 0 3 0 3 0 3
1 3
2 3 3
12 3 3 1 3 3 1 3 1 0 3 3 3
6 3 1 3 0 1 3
8 3 0 3 0 3 3 0 2
6 3 3 1 2 1 3
7 3 3 3 2 0 0 3
4 3 0 2 3
5 3 3 1 3 0
4 3 0 2 3
3 3 1 3
2 3 3
25 3 3 0 1 0 1 3 3 1 0 1 3 3 0 3 1 2 1 1 1 1 1 3 1 3
16 3 1 3 0 2 0 3 1 0 1 3 3 1 2 3 0
19 3 0 3 1 2 1 2 0 3 0 1 3 3 0 1 3 3 0 3
4 3 2 0 3
9 3 1 3 3 2 3 1 1 0
20 3 1 1 3 0 2 1 0 3 2 0 3 0 2 3 1 3 3 1 3
6 3 0 3 3 2 0
4 3 0 2 3
7 3 2 0 1 3 1 2
2 3 3
3 3 3 0
1 3
4 3 0 2 3
11 3 0 3 1 3 0 3 0 1 0 2
6 3 2 1 2 3 0
2 3 0
2 3 3
3 3 1 3
6 3 3 1 3 3 3
4 3 3 1 3
6 3 3 2 3 1 2
3 3 0 3
5 3 0 3 0 0
9 3 0 3 0 1 3 3 0 3
9 3 1 1 3 0 3 1 2 3
3 3 0 3
6 3 0 3 3 3 0
15 3 0 3 1 0 1 0 1 3 3 0 2 0 1 3
10 3 0 1 0 1 3 0 0 1 3
4 3 3 0 3
6 3 1 2 0 0 3
3 3 0 3
33 3 0 3 0 1 2 0 3 0 1 2 0 2 1 3 0 2 0 3 0 3 3 1 3 3 3 1 3 0 3 3 3 3
2 3 3
1 3
6 3 3 1 0 2 0
19 3 1 3 0 0 0 3 3 3 3 0 2 1 2 3 0 0 1 3
11 3 0 3 1 0 1 0 1 3 3 3
10 3 0 3 1 3 3 1 2 3 0
25 3 3 0 1 2 3 1 0 1 0 3 1 2 3 1 3 3 0 3 1 2 1 0 3 0
6 3 0 3 1 2 3
3 3 3 2
8 3 0 3 0 3 3 0 0
19 3 0 3 3 0 1 2 1 3 0 0 0 0 3 2 2 0 2 3
17 3 3 0 0 1 3 0 1 1 3 3 3 3 0 2 3 0
13 3 1 1 1 1 3 1 3 1 1 2 3 0
15 3 0 3 0 1 0 2 1 2 3 3 1 0 3 1
9 3 3 1 3 3 1 2 0 3
2 3 3
4 3 1 3 0
14 3 0 3 3 0 2 1 0 1 3 0 1 2 0
8 3 0 3 2 3 0 3 3
3 3 3 0
1 3
3 3 1 3
14 3 3 1 0 3 3 3 3 0 3 1 3 3 1
20 3 0 3 0 2 0 2 0 3 3 1 3 3 0 3 0 3 0 3 3
33 3 1 2 3 1 2 3 3 0 2 0 3 1 2 0 3 0 1 1 1 2 0 3 0 2 3 3 3 1 3 3 3 0
8 3 0 3 0 3 1 2 3
3 3 0 3
1 3
2 3 3
1 3
6 3 0 2 1 0 2
31 3 3 1 2 2 0 3 1 1 3 3 0 1 1 1 3 1 1 0 3 3 1 1 1 3 0 3 3 3 3 2
21 3 0 3 0 3 0 3 0 1 2 0 2 0 2 0 2 3 2 2 0 3
5 3 0 3 1 2
4 3 3 3 0
25 3 0 1 0 0 3 0 2 1 1 3 0 2 0 3 1 1 1 3 0 2 3 1 3 3
4 3 1 1 1
5 3 0 1 0 0
3 3 0 1
6 3 0 3 0 3 3
4 3 3 1 3
6 3 0 2 3 3 3
2 3 3
1 3
3 3 3 3
2 3 3
12 3 3 2 1 0 0 0 3 3 3 1 3
6 3 1 3 0 2 3
2 3 3
21 3 1 0 0 1 1 2 0 3 0 2 0 3 0 1 3 3 1 0 3 3
7 3 0 3 0 3 3 0
1 3
13 3 2 0 3 0 0 0 3 3 3 0 1 0
4 3 0 3 3
6 3 0 3 0 0 3
5 3 0 3 3 1
18 3 1 1 3 0 1 1 1 1 2 0 0 3 1 2 2 0 3
10 3 3 0 2 0 3 0 1 0 0
6 3 0 3 1 0 2
7 3 3 0 0 3 0 0
2 3 3
21 3 0 3 0 1 2 2 3 1 3 3 3 0 2 3 1 2 3 3 3 2
5 3 0 3 1 2
17 3 0 2 2 3 0 3 0 1 2 1 1 1 0 2 0 3
12 3 3 2 3 1 3 3 3 2 1 3 3
3 3 3 0
17 3 0 2 3 1 1 1 1 1 1 1 1 3 1 1 1 3
5 3 0 1 3 3
10 3 3 0 1 2 3 0 0 1 3
32 3 3 0 2 2 3 1 2 0 3 0 1 1 3 1 3 0 0 1 3 3 3 1 2 0 3 0 0 1 3 0 2
15 3 1 3 0 2 0 3 3 1 3 3 0 1 0 3
3 3 0 3
14 3 3 0 2 1 1 3 0 1 0 1 1 1 1
26 3 0 3 0 3 3 1 3 3 1 1 1 1 2 0 2 0 3 0 3 0 1 3 3 1 3
7 3 0 3 0 1 3 3
5 3 0 3 1 0
3 3 3 0
4 3 0 3 0
2 3 0
2 3 3
7 3 3 1 3 0 0 3
1 3
7 3 3 1 3 3 1 0
4 3 0 3 3
16 3 3 0 1 1 2 0 3 0 3 0 2 0 3 3 0
3 3 1 3
1 3
2 3 3
11 3 3 1 3 3 0 1 3 3 1 3
12 3 0 3 1 3 3 1 3 3 1 2 3
15 3 0 3 1 2 3 1 2 1 1 3 0 0 0 1
26 3 1 3 0 1 3 1 2 1 3 3 3 3 3 3 0 1 3 3 3 3 0 2 3 0 0
12 3 2 2 2 3 0 1 3 3 0 3 0
11 3 3 0 2 1 2 0 0 0 0 3
6 3 0 3 1 3 3
4 3 1 3 0
2 3 3
20 3 0 2 0 0 0 3 3 0 2 2 0 1 3 1 3 0 0 1 3
3 3 1 2
10 3 2 0 3 0 1 2 0 2 3
14 3 3 0 0 0 1 1 0 1 3 3 0 2 3
5 3 3 0 2 3
6 3 0 3 1 0 2
5 3 0 3 3 0
2 3 3
5 3 1 3 1 3
2 3 0
2 3 3
4 3 0 2 3
14 3 0 3 1 2 1 3 1 3 3 1 1 1 1
3 3 0 3
4 3 1 1 3
24 3 0 3 1 1 3 0 1 2 0 3 3 3 1 3 0 0 1 1 3 0 1 1 1
4 3 1 3 0
13 3 3 0 2 0 3 0 1 2 3 3 2 0
1 3
3 3 1 1
5 3 3 3 3 2
60 3 1 3 0 2 0 3 3 1 3 3 1 2 0 3 0 0 1 3 0 2 0 3 0 1 3 3 1 2 2 0 3 1 3 1 1 3 3 2 0 1 3 0 2 0 1 0 3 3 3 3 3 0 0 1 3 3 0 2 3
1 3
2 3 3
2 3 0
16 3 0 2 3 3 3 3 0 1 2 1 1 3 2 0 3
4 3 0 3 3
5 3 0 3 0 3
6 3 3 0 1 0 1
2 3 3
15 3 0 3 0 1 3 3 3 1 2 1 1 2 0 1
1 3
4 3 0 2 3
8 3 3 0 0 0 3 0 0
12 3 3 0 1 1 3 1 1 2 1 1 0
9 3 1 1 2 0 1 2 1 3
3 3 0 3
4 3 3 3 0
5 3 3 1 2 3
10 3 0 3 0 1 0 2 3 0 3
1 3
24 3 3 1 0 1 3 3 1 1 3 3 0 1 3 3 1 3 0 1 1 3 0 1 1
2 3 3
3 3 0 3
5 3 0 3 0 3
18 3 0 2 3 1 3 3 0 1 2 3 0 0 0 3 1 0 3
7 3 2 0 1 3 0 0
6 3 0 3 0 2 3
6 3 3 1 3 1 3
6 3 3 0 1 3 1
2 3 3
3 3 3 0
7 3 3 0 0 1 1 3
4 3 0 3 0
8 3 0 3 0 3 0 0 3
12 3 0 1 3 3 1 3 0 2 3 2 0
2 3 3
9 3 3 1 3 3 3 0 0 0
4 3 3 3 0
7 3 0 3 1 2 3 0
11 3 0 3 3 1 2 0 2 0 3 0
4 3 3 3 3
8 3 0 3 0 0 3 0 2
1 3
6 3 0 3 0 2 3
9 3 3 1 3 3 3 2 1 0
28 3 1 1 1 3 0 1 2 3 1 3 3 1 3 0 1 2 0 3 0 1 3 3 3 2 0 0 2
5 3 2 0 3 0
11 3 1 1 3 1 1 3 0 3 0 1
2 3 3
2 3 3
1 3
21 3 0 3 3 1 3 3 1 2 1 1 0 0 1 0 0 1 1 0 2 3
5 3 3 1 3 3
4 3 0 3 0
4 3 0 2 3
1 3
2 3 0
3 3 1 3
2 3 0
2 3 3
9 3 3 1 3 2 0 1 3 0
2 3 3
2 3 0
9 3 0 3 0 2 0 1 1 3
26 3 0 2 3 1 1 1 2 1 1 1 1 3 0 2 3 1 3 3 3 0 3 1 1 3 1
8 3 0 1 3 1 2 0 3
8 3 0 3 1 3 0 3 3
5 3 3 3 2 0
4 3 1 1 1
2 3 3
29 3 3 0 0 0 3 3 3 1 1 3 0 1 2 1 3 0 1 1 2 0 3 0 1 3 3 0 3 3
6 3 0 3 0 2 0
1 3
1 3
7 3 1 3 0 0 1 3
5 3 0 3 1 0
8 3 3 0 0 1 3 0 0
2 3 3
22 3 0 3 3 3 3 0 1 1 1 1 2 0 3 1 3 3 1 3 1 0 0
3 3 3 3
6 3 3 1 3 1 3
3 3 0 3
5 3 0 2 3 0
7 3 0 3 1 2 0 3
4 3 3 2 3
1 3
6 3 0 3 1 3 0
3 3 1 3
7 3 0 3 0 1 3 3
2 3 2
7 3 1 3 0 0 0 1
3 3 1 3
3 3 3 0
7 3 0 3 0 2 1 0
11 3 2 3 0 2 0 3 0 0 1 3
5 3 0 3 0 3
1 3
12 3 0 3 1 1 3 1 3 0 0 1 3
9 3 1 1 3 3 3 3 3 3
2 3 0
16 3 2 3 1 3 0 3 1 2 1 2 0 0 0 1 0
3 3 0 3
11 3 0 3 0 2 0 1 3 1 0 0
4 3 3 3 1
8 3 0 0 0 2 1 1 2
4 3 3 0 2
5 3 0 3 0 3
15 3 1 3 0 0 3 3 3 3 3 0 3 1 3 3
8 3 0 3 0 2 0 3 0
1 3
2 3 3
3 3 0 3
8 3 3 1 3 3 0 2 0
10 3 0 3 0 2 1 1 2 0 3
4 3 2 0 3
4 3 2 0 3
5 3 0 3 0 3
26 3 0 1 1 3 3 3 1 1 3 0 3 3 3 0 1 3 3 0 3 0 1 3 3 0 2
9 3 0 3 0 3 0 1 0 0
12 3 3 2 0 2 0 3 1 3 3 1 2
2 3 3
5 3 2 0 3 1
14 3 0 1 3 3 0 1 2 0 3 0 1 3 3
3 3 1 3
3 3 3 3
7 3 3 0 2 1 3 3
5 3 0 3 0 3
18 3 3 2 1 1 2 2 0 3 1 0 2 0 0 1 0 2 3
6 3 0 3 1 0 2
10 3 1 3 0 2 0 3 0 0 2
6 3 1 2 0 0 3
3 3 0 3
4 3 0 2 3
8 3 0 3 3 1 3 3 2
14 3 0 1 0 1 1 3 0 2 1 1 3 0 3
5 3 0 3 1 3
11 3 0 3 0 1 3 3 0 1 3 3
4 3 3 2 0
2 3 3
14 3 1 3 0 1 2 0 3 0 1 1 3 3 3
5 3 0 2 3 0
2 3 3
8 3 0 3 0 1 3 3 3
4 3 3 2 0
7 3 3 0 2 1 2 0
20 3 3 0 1 1 2 0 3 1 2 1 1 1 1 3 1 3 3 3 3
17 3 0 3 1 3 0 2 0 1 1 2 0 3 0 3 2 0
19 3 3 1 3 1 1 1 3 0 1 1 3 0 3 1 2 1 3 0
2 3 3
19 3 3 0 2 0 3 1 2 0 3 1 3 3 0 3 0 2 1 3
21 3 0 3 1 3 3 1 2 3 3 0 1 2 0 3 0 3 0 3 0 1
4 3 3 0 2
9 3 0 3 1 3 3 1 1 0
31 3 1 3 1 3 3 0 3 3 3 3 1 3 3 0 3 0 3 0 1 3 3 3 0 1 2 0 3 0 3 3
16 3 1 1 3 0 0 1 3 0 1 1 1 3 2 0 3
5 3 1 3 0 1
11 3 1 3 0 0 1 3 0 2 3 1
1 3
6 3 0 3 1 2 3
9 3 0 3 0 1 3 3 0 3
4 3 1 3 0
8 3 1 1 1 1 1 1 0
2 3 3
6 3 0 3 0 0 3
2 3 0
8 3 0 2 3 0 3 0 2
1 3
5 3 0 3 3 2
3 3 0 2
7 3 3 1 3 3 1 3
6 3 0 3 1 2 3
3 3 0 3
15 3 1 3 0 0 1 3 0 1 3 3 3 3 1 3
7 3 0 3 1 1 1 3
5 3 3 0 0 0
2 3 0
4 3 0 2 3
7 3 0 3 1 3 3 2
2 3 3
1 3
3 3 1 2
12 3 0 3 0 3 1 0 2 1 2 0 2
3 3 0 3
10 3 0 3 0 2 2 2 3 0 0
2 3 0
3 3 3 3
14 3 0 3 1 2 1 1 1 1 1 1 1 1 0
12 3 1 1 2 3 1 0 3 3 1 2 3
2 3 3
3 3 3 0
15 3 0 3 3 3 0 1 0 2 3 1 2 3 1 1
6 3 0 1 2 3 3
13 3 3 1 3 3 1 3 3 0 3 0 3 0
12 3 3 0 2 2 0 3 0 0 1 3 0
7 3 3 0 1 3 3 3
2 3 3
13 3 3 0 2 3 3 1 3 3 3 1 0 0
15 3 3 1 3 3 3 0 1 3 3 3 1 3 3 3
1 3
13 3 3 0 2 1 0 3 2 3 3 0 3 0
3 3 0 1
19 3 0 2 3 0 1 1 0 2 1 1 1 1 3 1 3 1 3 3
16 3 0 3 1 3 3 1 3 3 0 3 0 2 3 1 3
4 3 2 0 3
4 3 1 2 0
15 3 1 3 1 3 3 0 1 3 3 0 1 3 3 0
13 3 0 3 1 2 1 2 0 2 3 0 0 0
6 3 0 3 1 0 2
5 3 3 0 0 3
6 3 3 0 2 0 1
8 3 0 3 0 3 1 2 1
5 3 0 2 3 0
12 3 0 1 0 1 3 3 0 3 1 2 3
13 3 0 3 0 1 3 1 0 1 3 1 0 3
2 3 3
12 3 0 2 1 1 3 0 2 1 0 2 1
6 3 0 3 1 2 3
21 3 3 3 1 3 3 1 3 3 0 3 0 3 0 3 3 3 1 3 1 3
1 3
7 3 3 0 1 2 2 3
2 3 3
1 3
13 3 0 3 1 1 1 1 1 1 1 1 1 1
9 3 0 3 0 3 3 3 0 3
7 3 3 0 2 1 3 0
3 3 3 2
4 3 3 1 0
16 3 0 3 0 3 0 2 0 1 3 3 0 1 3 3 3
10 3 3 1 2 1 2 0 1 2 1
2 3 3
5 3 0 3 1 0
38 3 3 0 0 3 3 0 1 1 3 1 1 3 3 0 1 0 2 3 0 1 3 3 3 0 1 1 1 1 3 3 3 3 0 1 1 3 2
15 3 3 2 3 3 3 1 3 3 1 0 2 0 0 2
15 3 3 0 2 1 1 3 3 0 1 3 3 2 0 3
5 3 0 3 1 2
16 3 0 2 3 3 1 3 3 1 0 3 3 0 3 3 3
2 3 0
8 3 3 1 3 3 0 3 0
11 3 1 3 0 0 0 3 3 3 1 3
13 3 0 3 1 2 2 0 3 3 0 2 0 3
3 3 1 3
4 3 3 3 0
1 3
3 3 1 3
10 3 1 3 0 1 2 0 3 0 2
1 3
12 3 0 3 0 2 3 1 1 1 1 3 0
4 3 0 3 0
2 3 3
16 3 1 3 0 1 1 2 0 3 3 3 0 0 3 1 0
11 3 0 3 0 1 3 3 3 1 3 3
2 3 3
17 3 1 3 0 0 0 3 3 3 1 2 2 3 3 1 0 3
12 3 3 0 1 1 1 2 0 3 1 3 0
31 3 3 2 3 1 3 3 0 3 1 2 1 1 1 3 1 1 0 1 3 3 0 1 0 1 2 2 3 1 3 3
6 3 3 1 3 2 3
4 3 0 3 3
8 3 0 3 1 2 3 1 1
12 3 3 0 3 1 1 3 1 2 0 2 3
6 3 1 1 3 1 1
6 3 0 3 3 3 0
14 3 0 3 0 3 0 3 0 1 2 3 0 0 0
8 3 3 0 1 3 3 3 3
2 3 3
26 3 3 0 1 1 1 2 3 1 3 3 0 3 0 1 3 3 0 1 3 3 0 1 0 1 3
6 3 0 3 1 3 0
4 3 0 3 2
2 3 3
6 3 0 3 1 2 3
4 3 0 3 0
2 3 3
3 3 0 3
6 3 0 3 0 2 3
6 3 2 0 1 3 0
13 3 1 3 0 2 0 0 1 2 0 3 1 3
3 3 3 0
7 3 0 3 0 2 3 0
3 3 0 3
14 3 0 3 0 1 3 3 1 3 1 3 3 0 3
23 3 1 1 3 1 3 0 2 1 1 1 3 3 3 0 3 1 1 1 3 1 3 0
3 3 3 1
6 3 0 3 3 2 0
5 3 2 0 3 0
2 3 0
15 3 3 3 3 0 3 3 3 0 3 3 3 0 1 1
9 3 0 3 1 2 0 1 3 0
20 3 3 0 1 1 3 3 0 0 1 3 3 3 3 0 1 0 0 0 2
13 3 0 3 0 3 1 2 1 1 1 1 1 2
11 3 3 1 1 1 1 2 2 1 1 3
9 3 0 3 0 3 0 3 3 3
2 3 3
2 3 3
2 3 0
3 3 3 0
11 3 0 3 0 0 3 0 1 0 3 3
11 3 0 3 0 2 1 3 0 2 1 2
7 3 0 3 0 1 3 3
8 3 0 2 3 0 0 3 0
7 3 1 3 0 2 1 3
2 3 3
1 3
10 3 0 2 1 3 0 0 1 3 0
5 3 0 3 0 2
11 3 0 3 0 0 1 0 2 3 0 2
1 3
34 3 3 1 3 3 1 2 1 3 2 1 1 1 0 1 3 3 3 0 3 1 0 2 3 0 1 1 2 3 1 2 1 2 3
2 3 0
11 3 1 3 0 0 3 3 0 1 3 3
6 3 3 1 3 3 3
8 3 2 0 3 1 1 0 0
15 3 3 1 3 3 1 0 1 3 3 0 1 0 0 1
2 3 1
9 3 0 3 0 1 3 3 0 2
4 3 1 3 0
6 3 0 3 0 3 0
2 3 0
2 3 3
11 3 3 2 0 1 2 0 1 1 1 3
3 3 3 0
2 3 0
4 3 0 3 0
6 3 1 1 3 1 3
7 3 3 1 3 3 1 3
9 3 0 3 1 3 2 0 3 0
4 3 3 0 0
2 3 3
6 3 0 3 0 3 3
2 3 3
3 3 0 3
10 3 0 3 0 1 0 3 3 3 0
5 3 3 1 1 1
4 3 0 2 2
3 3 1 3
7 3 3 2 3 2 0 3
6 3 1 3 0 0 0
5 3 3 1 3 0
11 3 0 3 0 1 3 3 3 3 2 0
1 3
12 3 3 0 1 2 3 2 0 0 1 3 3
5 3 0 3 0 2
13 3 0 3 0 1 1 3 3 3 1 0 3 3
1 3
6 3 0 3 1 3 0
2 3 3
5 3 1 1 3 0
6 3 0 3 0 3 3
6 3 0 3 1 2 1
20 3 0 3 0 1 3 3 0 3 1 0 0 0 1 3 3 0 3 0 3
28 3 3 0 1 2 0 3 1 0 1 3 3 0 1 3 3 1 2 1 2 0 3 3 1 3 3 1 3
12 3 3 3 3 1 2 2 0 3 0 1 3
13 3 0 3 3 1 3 3 1 3 0 3 1 3
4 3 0 3 0
1 3
12 3 0 3 0 3 1 3 1 1 3 1 1
3 3 1 2
5 3 1 0 3 3
5 3 0 3 1 2
6 3 0 2 1 3 0
12 3 0 3 0 2 1 0 2 0 0 0 3
10 3 0 3 0 1 3 3 0 2 0
5 3 0 3 0 2
2 3 3
1 3
3 3 3 0
6 3 3 0 1 0 1
4 3 0 3 3
9 3 0 3 1 2 2 0 3 0
9 3 0 2 1 3 0 2 1 2
8 3 3 1 3 3 0 3 3
14 3 0 3 1 1 3 3 2 0 3 0 2 0 3
7 3 0 3 3 3 0 3
2 3 3
3 3 1 3
3 3 1 3
10 3 0 1 3 3 0 3 0 0 1
6 3 0 3 1 2 3
5 3 0 2 3 0
6 3 0 3 0 2 0
2 3 3
2 3 3
9 3 3 3 2 1 1 3 3 0
4 3 0 2 3
6 3 3 0 2 0 3
2 3 3
18 3 0 3 3 0 1 1 1 2 1 3 0 1 1 0 1 2 3
4 3 1 2 3
20 3 1 3 3 1 3 0 3 0 1 3 3 3 0 2 1 1 3 0 2
9 3 0 3 0 3 0 1 3 3
10 3 3 1 3 3 3 0 1 1 3
7 3 0 2 3 1 1 1
7 3 1 3 0 2 1 0
8 3 0 2 3 0 0 1 3
3 3 3 0
2 3 3
1 3
13 3 3 2 0 2 0 3 1 0 2 3 1 2
13 3 1 3 0 2 1 3 3 0 0 2 1 3
3 3 3 0
9 3 3 0 1 0 0 3 1 3
8 3 0 3 0 1 3 3 3
2 3 3
5 3 0 3 0 3
2 3 3
14 3 3 0 3 3 3 1 3 3 0 1 0 3 3
2 3 0
11 3 3 0 2 2 0 3 0 1 3 1
2 3 0
7 3 3 1 3 3 0 1
2 3 3
1 3
8 3 3 1 2 3 0 3 0
2 3 1
12 3 0 3 1 2 1 1 2 3 3 3 2
4 3 0 3 3
3 3 3 0
3 3 0 3
6 3 3 0 0 1 3
17 3 3 1 1 1 1 1 3 0 1 1 2 0 3 3 1 1
2 3 3
2 3 3
24 3 1 3 0 0 1 3 1 1 1 3 1 3 1 3 1 1 1 1 1 3 3 3 3
5 3 3 2 0 1
2 3 3
4 3 1 2 0
3 3 0 3
8 3 0 3 1 0 1 3 1
4 3 0 1 2
3 3 3 2
7 3 3 0 0 1 3 0
22 3 3 0 1 1 1 0 1 1 1 2 2 0 3 0 0 3 1 3 0 3 3
3 3 3 2
4 3 3 0 0
3 3 3 2
1 3
8 3 1 0 3 3 1 3 3
1 3
5 3 1 1 3 0
6 3 0 3 2 0 3
4 3 0 3 0
1 3
1 3
6 3 1 1 1 3 0
1 3
2 3 3
12 3 0 3 2 0 1 1 3 0 0 1 3
3 3 0 3
4 3 1 3 2
1 3
15 3 0 3 3 1 3 3 1 2 1 3 3 3 3 3
1 3
4 3 0 1 0
7 3 3 0 1 3 2 3
1 3
6 3 0 1 3 3 3
5 3 2 0 3 0
13 3 1 1 3 3 3 1 3 3 0 2 0 0
12 3 1 3 1 3 3 1 3 1 3 3 3
18 3 1 3 1 0 2 3 0 3 3 3 1 3 3 1 2 1 3
1 3
11 3 1 3 0 3 3 3 1 3 3 3
14 3 2 0 3 1 3 3 0 3 0 1 1 2 1
13 3 0 3 0 1 3 3 0 3 0 1 3 3
2 3 3
1 3
4 3 1 3 0
5 3 3 0 2 0
4 3 0 3 0
2 3 2
3 3 0 3
11 3 1 1 3 0 3 0 0 1 3 1
11 3 1 1 1 1 1 3 3 3 0 3
3 3 0 3
4 3 0 3 0
16 3 0 3 1 0 1 2 2 0 3 1 3 0 3 3 0
1 3
4 3 0 2 3
3 3 0 3
6 3 0 2 1 3 0
5 3 0 3 0 3
3 3 0 3
8 3 0 1 0 3 3 1 3
5 3 0 3 1 3
3 3 3 0
3 3 3 0
2 3 3
8 3 3 0 1 2 0 3 3
1 3
2 3 3
2 3 3
3 3 1 3
1 3
16 3 0 3 0 3 0 1 0 1 3 3 3 0 2 3 3
5 3 0 2 3 0
5 3 0 3 1 2
14 3 3 0 0 0 3 3 3 3 1 3 3 3 0
8 3 1 3 0 2 0 2 3
2 3 3
5 3 3 0 3 3
4 3 3 0 0
7 3 0 3 3 0 2 1
3 3 0 2
8 3 1 3 0 3 3 1 0
2 3 3
8 3 1 3 0 2 1 3 0
5 3 3 0 0 3
15 3 0 3 0 3 0 3 0 1 3 3 1 2 0 3
14 3 2 2 1 0 1 2 3 0 2 3 0 1 0
3 3 1 3
12 3 3 0 2 1 1 3 3 3 3 3 2
20 3 1 1 3 0 1 3 2 1 1 3 3 3 3 0 3 0 1 2 3
9 3 3 1 3 0 3 0 2 1
2 3 3
16 3 3 1 3 0 2 0 0 1 3 3 3 0 2 0 3
1 3
16 3 0 3 1 3 3 3 3 0 0 3 1 2 1 0 1
3 3 3 3
5 3 0 3 0 1
3 3 1 3
6 3 0 3 3 0 0
12 3 0 1 2 0 1 1 3 3 0 1 0
3 3 3 2
2 3 3
11 3 0 3 3 1 3 3 0 2 0 3
4 3 0 3 0
7 3 0 3 1 2 1 0
8 3 3 0 2 2 0 3 3
11 3 3 0 1 1 2 0 3 1 3 0
13 3 0 3 0 1 3 3 1 2 2 0 2 3
3 3 1 3
8 3 0 3 0 1 3 3 3
13 3 3 0 0 3 3 3 2 2 1 3 1 3
3 3 3 0
4 3 1 1 3
15 3 0 1 1 2 0 3 0 3 1 3 0 0 1 3
11 3 0 3 0 2 0 3 0 0 1 3
4 3 2 0 3
6 3 1 3 3 2 0
8 3 0 3 0 2 0 3 0
14 3 0 3 0 1 1 1 1 1 2 3 1 3 1
8 3 0 1 3 3 1 2 0
5 3 1 1 3 0
12 3 3 1 3 3 0 1 3 3 3 0 0
2 3 3
3 3 3 0
3 3 0 1
14 3 1 3 1 3 3 3 1 2 3 0 0 1 3
12 3 3 1 0 1 1 2 3 0 0 0 2
44 3 0 3 0 1 3 3 1 1 0 3 0 0 1 3 3 3 3 0 1 1 2 3 1 1 3 0 1 3 3 0 3 0 0 3 1 3 0 3 3 1 3 3 3
4 3 1 1 3
8 3 0 3 1 0 1 3 3
3 3 1 3
9 3 3 1 3 0 3 0 1 2
2 3 3
2 3 3
2 3 3
5 3 1 3 0 0
6 3 3 0 2 0 1
5 3 0 3 0 3
4 3 1 1 3
20 3 1 3 0 1 0 1 3 1 3 0 2 1 0 2 2 1 3 0 0
3 3 3 3
5 3 1 1 3 3
4 3 1 2 0
15 3 3 0 2 0 3 0 0 3 0 1 0 1 0 2
1 3
1 3
5 3 0 3 3 3
4 3 0 2 3
1 3
2 3 3
11 3 0 3 1 3 3 0 0 1 3 0
12 3 1 3 0 2 0 2 3 0 3 3 0
16 3 3 0 0 1 1 3 1 3 3 3 1 3 2 2 0
5 3 3 0 1 1
9 3 3 0 1 1 1 1 2 3
4 3 0 2 3
7 3 0 3 0 3 3 0
10 3 0 3 1 3 1 2 0 1 0
4 3 3 2 3
5 3 1 1 3 0
3 3 0 1
2 3 1
2 3 3
11 3 0 3 3 0 1 2 0 2 3 0
2 3 1
3 3 3 0
3 3 0 3
18 3 0 3 3 3 0 3 0 1 3 3 0 1 0 0 2 0 3
4 3 0 3 0
2 3 3
9 3 3 1 2 0 3 0 1 0
6 3 3 0 0 3 0
8 3 0 3 0 1 3 3 3
6 3 0 3 1 2 3
4 3 1 0 0
3 3 0 3
3 3 3 0
11 3 0 2 0 1 2 2 0 3 3 3
3 3 3 0
9 3 1 3 0 2 3 1 0 3
4 3 0 2 3
19 3 3 0 0 3 3 0 0 3 0 2 1 0 2 0 0 1 0 0
7 3 3 0 0 3 3 3
12 3 0 2 3 0 0 3 0 0 2 0 1
13 3 0 3 0 2 3 1 2 0 1 1 1 3
3 3 3 2
3 3 3 0
4 3 0 3 3
1 3
16 3 0 2 3 3 3 3 1 3 0 1 2 0 2 2 1
12 3 0 2 1 1 3 0 2 0 1 3 3
5 3 1 1 3 0
2 3 3
2 3 3
2 3 3
5 3 3 0 0 0
6 3 3 0 2 2 0
10 3 0 3 3 3 0 0 1 3 0
7 3 0 2 3 1 0 3
18 3 1 1 3 1 3 3 0 3 1 0 1 3 3 1 2 3 0
3 3 0 1
7 3 3 1 3 3 1 3
3 3 0 3
27 3 0 3 0 1 2 2 0 3 0 1 0 3 3 1 3 0 3 0 3 0 1 3 3 0 0 3
17 3 2 0 1 3 0 1 2 3 2 3 0 1 2 3 0 0
15 3 0 3 0 1 2 0 2 3 1 1 3 0 2 3
9 3 3 1 3 0 1 2 0 2
3 3 1 3
1 3
8 3 1 2 0 2 2 0 3
10 3 3 1 3 3 0 3 0 3 3
2 3 3
1 3
4 3 1 1 3
2 3 3
8 3 2 0 3 0 0 1 3
10 3 0 3 1 2 1 2 2 3 0
8 3 0 3 1 0 1 0 2
5 3 0 2 0 2
8 3 1 3 0 1 2 3 0
2 3 3
31 3 0 3 1 3 0 0 2 3 0 2 0 3 1 2 1 3 0 1 1 1 1 0 1 1 0 0 3 0 1 2
12 3 0 3 1 2 1 1 0 3 3 0 3
25 3 3 1 1 3 0 3 3 3 3 0 1 1 1 2 3 0 1 1 3 3 2 0 0 3
1 3
7 3 0 3 1 3 1 3
1 3
8 3 3 1 3 1 0 2 0
2 3 3
6 3 3 0 0 1 3
29 3 0 3 1 3 1 2 0 1 1 2 0 3 0 1 2 0 2 0 3 1 2 1 1 2 0 3 3 2
3 3 3 0
2 3 0
5 3 0 3 0 2
37 3 1 3 0 0 3 3 0 1 3 2 3 0 1 3 0 0 1 3 0 0 3 3 0 3 0 2 3 2 0 0 1 2 2 0 1 1
23 3 0 2 1 3 0 2 0 3 0 3 3 1 3 3 0 2 0 3 1 2 2 0
11 3 1 3 1 3 3 3 0 2 0 3
1 3
3 3 1 3
3 3 3 3
2 3 0
6 3 1 1 3 3 0
2 3 0
10 3 0 3 1 2 0 3 0 0 0
5 3 0 2 3 0
8 3 0 3 1 3 0 2 3
3 3 1 3
3 3 3 0
4 3 3 2 0
2 3 3
5 3 0 2 3 0
3 3 3 0
11 3 3 1 2 1 1 1 2 0 3 0
4 3 3 0 2
27 3 0 3 0 2 0 3 0 1 1 1 0 1 2 3 1 3 3 0 1 3 3 1 3 0 0 0
2 3 0
4 3 0 3 3
4 3 0 3 0
1 3
2 3 3
5 3 3 1 3 3
7 3 0 3 3 0 2 0
9 3 3 1 3 3 1 3 1 3
3 3 3 0
1 3
3 3 1 3
13 3 3 1 3 3 3 2 1 3 3 0 3 0
13 3 0 3 0 3 0 3 0 1 2 1 0 3
3 3 0 3
18 3 0 0 2 3 0 0 1 3 0 1 1 3 1 0 1 0 3
13 3 0 3 0 1 3 3 0 0 2 3 1 1
3 3 3 0
3 3 0 3
4 3 0 3 3
4 3 1 3 0
12 3 0 3 0 1 2 2 1 3 0 0 0
12 3 3 0 2 2 0 0 3 1 3 3 0
15 3 0 3 0 1 3 3 1 2 1 3 2 0 2 3
2 3 3
6 3 0 3 1 3 3
11 3 0 3 0 2 0 3 0 1 2 3
1 3
7 3 2 0 3 0 2 1
2 3 3
3 3 0 3
3 3 0 3
11 3 0 3 0 2 3 0 1 3 3 3
8 3 3 1 3 3 1 3 0
2 3 3
12 3 1 1 0 3 0 0 1 2 1 1 3
3 3 0 3
3 3 3 0
4 3 3 2 3
3 3 0 3
18 3 3 3 0 1 1 2 0 3 3 0 1 2 3 1 3 3 3
12 3 0 3 1 0 1 3 1 0 1 3 0
6 3 3 0 0 3 3
6 3 0 3 0 2 1
32 3 0 3 3 0 1 1 1 1 1 1 3 3 3 3 0 3 1 2 0 3 0 2 0 3 1 0 2 3 2 0 3
2 3 3
15 3 0 2 3 3 1 1 3 0 2 0 3 3 2 1
2 3 3
3 3 3 0
12 3 3 1 0 2 0 1 3 3 0 2 3
2 3 3
2 3 3
2 3 3
1 3
36 3 3 0 1 0 2 0 3 0 1 3 3 0 1 3 3 1 3 1 1 3 3 2 1 1 3 2 1 1 1 1 1 3 1 3 0
7 3 1 1 1 1 0 0
12 3 0 1 1 3 3 3 0 3 0 1 2
2 3 3
3 3 3 0
2 3 3
9 3 0 3 1 0 1 0 3 2
11 3 0 2 3 1 3 3 2 0 3 0
7 3 3 1 3 3 1 3
5 3 1 3 0 2
12 3 1 1 1 3 0 3 0 1 3 3 0
27 3 0 3 1 3 1 0 2 0 0 3 3 3 3 0 3 3 2 0 1 3 0 0 3 0 0 3
5 3 0 3 0 0
11 3 0 3 1 3 0 3 0 1 3 3
6 3 0 2 1 1 3
3 3 3 0
2 3 3
11 3 3 1 3 0 2 1 3 0 2 0
4 3 1 1 3
9 3 0 3 1 3 0 3 3 2
18 3 3 1 3 3 1 1 3 0 2 0 3 1 0 1 0 0 1
2 3 1
8 3 0 3 0 1 2 3 3
1 3
23 3 3 1 3 3 0 3 0 3 0 3 2 3 1 3 3 1 1 1 0 1 2 3
7 3 3 0 1 3 2 3
4 3 1 1 3
27 3 3 1 3 3 3 1 3 3 0 3 0 3 1 0 1 3 3 0 3 0 0 3 0 2 0 3
2 3 3
4 3 3 0 2
5 3 3 0 0 0
7 3 0 3 0 3 0 2
2 3 3
14 3 0 3 1 2 1 2 3 2 0 1 3 0 3
2 3 2
8 3 3 1 3 3 1 2 3
10 3 1 3 1 1 3 3 3 0 0
1 3
3 3 0 1
3 3 2 2
4 3 0 3 0
3 3 1 1
5 3 2 0 1 3
6 3 3 1 3 3 3
6 3 3 0 3 3 3
9 3 1 1 3 3 0 3 1 3
13 3 1 0 2 3 0 2 3 0 1 2 0 3
3 3 3 0
8 3 3 0 1 3 1 0 3
3 3 1 3
19 3 0 3 1 0 1 3 3 0 3 0 3 0 3 1 2 1 1 3
2 3 3
2 3 3
16 3 0 3 0 1 3 3 1 0 1 2 1 1 2 1 3
20 3 3 1 3 3 3 1 3 0 3 1 2 1 1 2 0 3 3 2 0
12 3 3 0 0 1 3 0 1 2 3 0 0
3 3 3 0
2 3 2
3 3 0 3
30 3 0 3 3 0 2 0 3 1 2 2 1 1 3 0 0 3 3 0 1 3 3 3 1 3 3 0 3 0 2
3 3 0 3
11 3 3 3 3 2 1 0 1 3 3 3
5 3 0 2 0 0
3 3 0 3
4 3 0 2 3
3 3 0 3
3 3 3 2
4 3 2 0 3
11 3 0 2 3 0 1 1 2 0 2 3
1 3
26 3 2 0 3 0 0 0 0 3 0 1 2 3 3 0 2 0 3 0 3 1 3 3 3 3 0
4 3 3 3 3
16 3 3 1 1 3 2 3 0 2 1 1 3 0 3 3 0
3 3 3 0
9 3 3 3 1 3 1 2 3 2
4 3 3 0 2
6 3 0 3 0 3 3
3 3 3 0
7 3 1 3 0 2 1 2
6 3 3 1 3 3 3
1 3
27 3 0 3 0 2 0 1 3 0 2 3 0 3 0 1 3 3 0 1 3 3 3 1 3 3 2 3
4 3 1 3 0
12 3 0 3 1 0 1 1 1 1 2 3 2
21 3 3 1 3 3 0 3 0 2 0 1 3 0 3 0 3 0 3 3 0 0
2 3 3
2 3 3
16 3 1 3 0 2 3 1 3 0 0 1 3 3 3 0 2
3 3 3 2
4 3 3 0 0
12 3 0 3 1 3 0 3 1 2 0 3 0
5 3 3 0 2 1
5 3 3 3 0 1
3 3 1 3
5 3 1 1 3 0
40 3 0 3 0 3 1 0 1 2 2 3 0 3 1 3 3 0 0 1 1 2 0 1 2 1 1 3 3 3 3 0 3 2 0 3 0 1 1 0 2
3 3 3 2
2 3 3
13 3 3 3 1 3 3 0 1 3 3 1 3 3
4 3 3 0 2
2 3 0
6 3 2 0 3 1 1
21 3 3 2 3 1 1 3 3 0 3 3 0 2 2 0 0 3 1 3 3 0
22 3 0 2 3 0 1 1 2 3 0 0 3 3 1 2 0 1 3 0 0 3 0
2 3 3
4 3 1 3 0
8 3 0 3 1 3 0 2 3
5 3 1 3 0 2
6 3 0 3 1 3 0
1 3
10 3 1 3 0 2 0 1 2 3 1
1 3
5 3 0 3 0 3
14 3 0 3 0 1 3 3 0 3 1 0 1 3 3
3 3 3 1
2 3 1
2 3 3
12 3 0 3 1 0 1 0 1 3 3 0 3
3 3 0 3
11 3 3 0 2 0 3 1 3 0 2 3
7 3 3 2 0 0 2 2
4 3 0 1 2
15 3 3 0 3 1 1 1 1 1 1 3 1 3 0 0
12 3 1 3 1 3 3 0 1 3 3 0 3
7 3 1 3 1 3 1 3
32 3 0 2 3 0 1 3 1 3 3 3 1 3 0 3 0 1 2 3 1 2 0 1 1 1 1 2 0 3 0 2 3
2 3 3
6 3 1 1 3 3 2
9 3 0 3 0 1 2 0 1 1
6 3 0 1 0 1 3
1 3
6 3 0 3 2 0 3
10 3 1 3 0 2 2 0 3 0 0
4 3 3 1 2
3 3 0 3
12 3 0 1 3 3 1 2 1 2 1 3 0
10 3 0 3 1 0 1 3 3 3 0
3 3 1 3
1 3
7 3 1 3 0 2 0 3
6 3 2 0 1 3 0
1 3
2 3 3
11 3 0 3 1 3 0 2 1 3 0 2
19 3 0 0 2 2 3 1 3 1 3 0 0 3 3 0 1 3 0 0
12 3 3 0 3 3 3 0 2 3 1 3 3
15 3 0 2 3 0 1 1 1 2 0 3 0 3 0 2
3 3 3 2
19 3 3 0 1 3 3 1 1 1 1 1 3 2 1 0 1 3 3 3
2 3 0
1 3
6 3 0 3 1 2 3
5 3 0 3 1 3
15 3 3 0 2 3 1 0 3 0 1 2 1 3 0 2
10 3 3 0 1 2 0 3 0 3 0
15 3 0 3 3 0 1 1 1 1 3 2 1 1 3 1
2 3 3
4 3 3 1 3
6 3 1 1 3 3 0
5 3 3 0 0 3
18 3 0 3 1 3 3 2 0 1 1 1 1 1 0 1 0 3 2
8 3 1 3 0 0 3 3 3
21 3 0 3 1 2 1 3 0 1 2 0 3 0 2 3 3 0 1 2 3 0
2 3 3
18 3 3 0 1 3 2 1 3 1 3 3 0 3 0 1 3 3 3
1 3
7 3 1 1 1 3 2 3
10 3 3 0 1 0 1 1 2 0 3
4 3 3 0 1
3 3 0 3
4 3 3 0 0
3 3 0 3
1 3
3 3 1 3
30 3 0 3 0 3 0 1 1 1 1 3 3 0 1 2 0 3 0 0 0 3 3 3 0 3 0 2 3 0 3
11 3 3 0 0 0 3 3 3 2 0 3
6 3 1 3 0 0 0
3 3 0 3
3 3 1 3
2 3 3
15 3 0 3 0 1 2 0 3 1 1 3 3 0 2 0
3 3 1 3
20 3 3 0 2 0 3 1 3 0 1 0 1 1 0 1 3 3 1 1 3
4 3 0 2 3
22 3 3 0 0 1 3 1 3 3 1 1 3 3 1 2 2 0 3 1 2 1 0
8 3 3 0 0 0 1 0 3
2 3 3
4 3 3 0 2
11 3 0 3 0 2 3 1 1 3 3 3
11 3 3 0 0 3 3 1 0 2 1 0
5 3 0 3 0 2
4 3 1 1 3
2 3 3
4 3 3 0 2
4 3 1 1 3
2 3 3
2 3 3
19 3 0 2 3 0 1 1 1 1 1 0 2 1 3 1 3 3 0 3
15 3 3 1 3 3 0 3 1 3 1 1 3 0 3 3
1 3
6 3 0 3 1 3 0
15 3 0 1 1 1 0 2 0 3 1 2 2 0 3 0
6 3 3 0 2 0 3
3 3 0 3
2 3 3
22 3 3 1 3 0 0 0 1 3 3 1 2 2 0 3 0 2 1 3 1 3 0
4 3 0 3 3
5 3 1 1 1 3
2 3 0
3 3 0 3
8 3 3 0 2 1 0 3 3
4 3 3 0 2
2 3 3
3 3 3 2
12 3 1 3 0 2 0 3 0 1 2 0 3
23 3 1 2 0 0 0 3 3 3 1 2 3 0 2 1 0 1 3 0 2 1 2 0
17 3 0 3 1 2 1 1 2 3 1 3 3 1 2 3 2 1
9 3 0 3 0 1 2 0 3 0
7 3 0 3 0 1 1 3
8 3 0 3 1 3 3 2 0
4 3 0 3 3
2 3 0
1 3
10 3 0 3 1 2 3 0 2 0 3
4 3 3 0 0
5 3 0 3 1 3
32 3 3 1 0 0 3 0 0 2 0 3 1 3 1 3 0 1 3 3 3 0 2 1 3 0 2 2 2 0 1 3 3
8 3 0 3 0 2 3 2 2
18 3 3 2 0 0 1 3 3 1 0 1 2 3 1 3 1 3 3
3 3 0 3
3 3 1 3
7 3 0 3 0 3 1 2
6 3 0 3 0 2 2
2 3 3
4 3 0 1 1
1 3
4 3 3 2 0
2 3 3
10 3 3 0 2 0 3 1 2 1 0
8 3 0 3 1 0 0 2 3
2 3 3
1 3
14 3 3 0 1 3 1 1 0 1 3 3 1 1 3
18 3 1 1 3 1 1 1 0 1 1 0 1 2 0 1 0 1 3
11 3 0 2 3 2 0 3 0 0 3 0
2 3 3
8 3 0 3 1 3 1 1 1
3 3 0 3
2 3 3
5 3 3 1 3 3
2 3 3
6 3 0 3 3 0 2
6 3 0 3 1 2 1
4 3 1 1 3
5 3 3 0 0 0
3 3 3 2
1 3
6 3 2 0 1 3 0
5 3 1 1 1 1
6 3 3 0 1 1 0
4 3 3 2 3
2 3 3
3 3 3 2
2 3 3
2 3 3
7 3 3 0 1 1 3 1
3 3 1 3
9 3 3 1 3 3 0 1 0 2
17 3 0 3 1 0 1 3 3 0 3 0 1 3 1 2 3 2
12 3 0 2 3 0 2 1 1 1 3 0 3
10 3 0 2 3 0 2 1 1 1 1
2 3 0
2 3 3
11 3 0 3 0 1 3 3 0 3 1 3
9 3 1 3 1 2 3 3 3 2
1 3
7 3 0 1 2 3 0 0
1 3
3 3 3 2
3 3 1 1
7 3 1 3 1 2 3 3
3 3 0 3
4 3 2 0 3
7 3 0 3 1 3 3 0
3 3 3 0
13 3 0 0 2 3 0 1 0 1 2 1 1 0
20 3 0 3 0 1 3 3 1 3 0 1 1 0 1 3 3 3 1 3 3
6 3 1 3 0 2 1
8 3 3 0 1 1 3 1 3
1 3
3 3 1 2
3 3 0 3
2 3 3
12 3 3 3 0 1 3 0 3 2 2 0 1
2 3 3
8 3 1 3 1 3 3 3 2
8 3 0 2 3 0 1 1 0
4 3 3 0 0
3 3 0 3
9 3 3 0 2 0 3 3 3 3
9 3 3 0 1 2 3 0 0 0
5 3 1 1 3 0
24 3 0 3 1 2 2 0 3 1 1 1 1 1 3 3 2 1 2 0 3 1 0 2 0
3 3 1 3
2 3 3
15 3 1 1 3 0 0 3 3 1 1 2 3 1 3 3
5 3 0 3 1 3
8 3 0 3 0 3 3 1 2
3 3 1 2
9 3 0 3 0 1 2 3 0 1
5 3 0 3 1 3
6 3 3 0 1 0 3
1 3
15 3 0 3 1 1 1 3 0 1 1 3 0 3 0 2
3 3 0 1
4 3 1 1 2
6 3 0 2 1 3 0
4 3 3 0 2
10 3 0 3 0 1 3 3 0 3 3
4 3 1 1 3
16 3 0 3 0 1 2 0 1 1 1 1 1 2 0 0 3
8 3 3 0 0 1 3 0 0
11 3 1 3 1 1 1 1 1 3 1 3
15 3 0 3 1 0 2 3 2 1 2 0 3 0 2 0
5 3 3 1 3 3
10 3 3 0 1 2 0 2 3 0 0
3 3 0 3
3 3 3 0
9 3 0 3 1 2 1 2 0 1
13 3 1 1 2 0 3 0 1 3 3 1 1 3
2 3 3
3 3 1 2
10 3 3 1 2 1 3 3 3 3 0
2 3 3
13 3 1 0 3 3 0 1 1 3 1 1 1 3
2 3 3
10 3 0 3 0 0 3 0 2 3 0
3 3 0 3
3 3 0 3
5 3 1 3 0 0
17 3 3 2 0 0 3 3 0 3 0 2 0 2 3 0 2 3
3 3 1 3
3 3 1 3
11 3 3 1 0 1 2 1 1 3 3 0
7 3 0 2 3 1 1 3
11 3 0 3 0 2 3 1 3 3 0 3
25 3 3 1 3 3 0 3 1 3 0 0 3 3 1 0 1 0 2 0 0 1 3 3 0 2
3 3 0 3
10 3 1 3 2 0 2 0 3 3 3
13 3 1 3 1 3 3 1 3 0 1 2 0 3
9 3 3 1 2 2 0 0 2 3
17 3 0 3 3 1 3 3 1 0 2 0 0 0 3 3 1 1
5 3 0 3 0 3
3 3 0 1
2 3 3
10 3 1 1 3 0 3 1 2 0 3
2 3 3
2 3 3
9 3 0 3 0 3 3 3 0 2
4 3 2 0 3
6 3 0 3 0 1 0
21 3 0 3 0 3 1 2 2 0 3 0 1 1 3 3 3 3 3 3 3 0
18 3 0 3 0 2 0 2 1 1 3 3 3 3 0 1 3 3 3
18 3 3 1 3 3 3 3 3 3 3 3 3 1 3 0 2 3 0
2 3 3
10 3 0 3 0 3 0 3 2 0 3
18 3 0 3 0 1 3 3 1 0 1 3 3 0 1 3 3 3 0
2 3 3
5 3 0 2 3 0
5 3 1 3 0 0
1 3
8 3 3 0 1 1 1 1 1
14 3 3 2 1 3 2 0 3 1 3 3 0 0 0
4 3 0 2 3
7 3 3 0 1 1 1 2
15 3 0 3 0 1 3 3 0 1 3 3 0 1 2 3
3 3 1 3
7 3 0 3 1 2 0 3
5 3 1 3 1 0
12 3 3 0 2 0 3 1 2 2 3 2 1
3 3 0 3
1 3
1 3
1 3
1 3
2 3 3
9 3 0 3 0 1 2 2 0 3
8 3 3 1 3 3 1 2 3
3 3 3 0
18 3 3 1 3 3 1 2 0 3 0 1 1 3 0 2 2 2 3
8 3 1 1 3 0 0 0 3
6 3 0 3 1 0 2
3 3 1 3
9 3 3 0 2 0 1 2 0 3
6 3 0 3 1 3 3
7 3 3 0 1 1 0 2
4 3 0 3 3
3 3 3 0
21 3 0 1 3 3 0 1 3 3 0 3 3 3 0 3 0 1 3 3 3 0
2 3 3
13 3 0 3 0 2 3 0 1 3 3 3 3 0
1 3
14 3 2 3 0 1 3 3 1 1 3 0 3 0 0
2 3 0
19 3 0 2 1 3 0 1 1 1 2 0 3 0 0 3 1 3 1 3
2 3 3
9 3 0 3 0 2 0 0 2 0
1 3
22 3 3 0 2 0 3 0 1 0 1 3 3 0 1 1 1 3 3 3 0 3 0
15 3 0 3 1 2 1 1 0 1 1 2 1 3 1 3
2 3 3
3 3 3 2
6 3 1 1 3 3 3
1 3
3 3 3 1
10 3 3 0 2 0 0 2 3 0 2
15 3 0 3 3 0 1 1 1 1 1 2 0 3 3 0
4 3 3 0 0
33 3 1 3 1 3 0 3 0 1 3 3 1 1 1 3 1 1 3 0 2 1 1 3 0 1 0 1 2 1 2 0 3 0
3 3 0 3
1 3
2 3 0
15 3 3 1 1 3 0 1 0 2 0 3 1 3 3 0
11 3 3 0 0 3 3 1 1 1 1 1
6 3 1 1 1 1 3
4 3 0 3 3
12 3 0 3 0 3 0 3 3 1 3 3 0
9 3 1 0 3 1 0 3 0 3
9 3 1 3 0 0 1 1 3 0
6 3 0 3 1 2 3
3 3 1 2
2 3 0
3 3 3 0
6 3 1 1 1 3 0
21 3 0 0 0 3 2 1 1 1 1 1 2 3 2 0 0 0 0 1 2 3
10 3 0 3 0 2 0 2 1 1 0
6 3 3 0 1 0 2
2 3 3
2 3 3
7 3 1 3 0 2 3 3
10 3 0 3 0 1 0 1 3 3 3
6 3 3 0 3 3 3
1 3
9 3 0 3 1 3 0 0 3 3
5 3 0 3 1 2
17 3 0 1 3 3 0 2 0 1 3 0 2 0 1 2 3 0
8 3 0 3 1 2 0 3 0
2 3 3
2 3 3
4 3 3 0 0
23 3 1 1 3 0 2 0 2 3 0 1 2 3 0 1 3 3 0 3 0 1 3 3
6 3 0 3 3 0 1
3 3 3 0
5 3 0 3 0 0
5 3 3 0 0 3
4 3 0 2 3
4 3 1 1 3
16 3 0 3 1 2 1 1 2 0 3 0 1 3 3 0 3
7 3 3 0 1 1 2 0
3 3 3 2
13 3 0 3 0 1 3 3 0 2 1 0 0 3
4 3 0 2 3
2 3 3
19 3 0 2 1 3 0 1 3 3 3 1 0 0 1 1 0 1 3 3
8 3 0 3 0 3 1 3 3
12 3 0 3 0 2 0 1 3 0 3 1 2
8 3 3 0 1 2 1 3 0
11 3 0 3 0 2 0 1 3 0 0 0
5 3 0 3 3 0
4 3 0 3 3
4 3 0 3 0
17 3 0 3 0 1 3 3 0 1 3 3 0 3 0 2 3 0
6 3 1 1 3 0 2
3 3 3 3
5 3 0 3 3 0
8 3 0 1 3 3 1 3 0
6 3 3 1 0 2 3
24 3 3 1 3 3 0 3 3 0 1 1 1 1 1 1 2 0 2 3 0 2 0 2 3
5 3 3 1 3 3
4 3 3 0 2
7 3 1 2 0 1 1 2
13 3 3 0 1 1 1 1 1 1 1 2 0 3
3 3 0 3
3 3 1 3
6 3 0 3 0 1 1
2 3 3
4 3 0 1 0
6 3 0 3 0 3 0
2 3 3
3 3 3 0
4 3 3 2 3
3 3 3 0
7 3 0 3 1 3 1 3
5 3 0 3 1 2
5 3 0 3 1 2
6 3 0 3 3 1 2
14 3 1 3 0 2 0 3 3 1 3 3 0 1 0
7 3 0 3 1 2 1 3
4 3 1 3 0
3 3 3 0
3 3 0 3
8 3 0 3 0 1 1 0 3
3 3 1 2
6 3 0 3 0 3 0
21 3 0 3 0 3 0 0 3 1 0 1 3 3 1 1 3 3 0 0 0 3
6 3 3 1 1 3 3
9 3 0 3 0 3 0 1 3 2
2 3 3
13 3 3 0 0 3 0 0 2 0 3 1 1 3
4 3 0 3 3
20 3 0 3 0 2 3 2 0 1 3 0 1 1 3 0 1 3 3 0 1
9 3 0 3 0 1 3 3 0 2
11 3 1 3 0 1 1 1 3 1 1 3
6 3 0 3 3 0 2
9 3 2 0 3 0 2 3 2 3
10 3 0 3 0 3 1 3 0 2 3
10 3 0 2 1 3 1 1 3 3 3
9 3 0 3 1 2 1 1 0 1
4 3 3 0 2
8 3 0 3 1 3 0 1 0
3 3 3 1
3 3 0 3
3 3 1 3
11 3 0 3 3 1 3 3 0 1 1 3
6 3 0 3 1 2 3
4 3 3 1 2
11 3 0 3 1 0 1 3 3 2 0 3
10 3 0 3 1 3 0 3 1 2 3
1 3
3 3 1 3
4 3 1 1 3
1 3
7 3 0 3 0 2 0 3
9 3 3 0 1 3 2 0 1 3
21 3 3 1 3 3 1 0 3 3 0 1 3 3 0 1 3 3 3 1 3 3
5 3 0 1 2 3
2 3 3
2 3 3
4 3 1 0 0
2 3 3
3 3 1 3
4 3 0 3 0
4 3 0 3 0
11 3 0 1 3 1 0 3 3 1 3 3
2 3 3
4 3 3 3 1
7 3 0 3 1 1 1 1
2 3 3
9 3 3 0 1 0 2 0 3 3
3 3 0 3
21 3 1 3 0 2 3 2 0 0 3 3 1 1 2 1 1 2 0 2 1 3
10 3 3 3 1 3 3 3 0 1 3
1 3
2 3 3
11 3 0 3 0 2 3 1 1 3 3 0
2 3 3
27 3 0 2 3 0 1 1 1 1 1 3 3 3 3 1 3 1 3 3 0 1 3 3 0 1 3 1
6 3 3 0 1 1 1
2 3 3
1 3
1 3
11 3 0 3 1 2 2 3 2 3 3 3
3 3 1 3
5 3 1 1 1 3
9 3 1 1 3 3 0 2 1 2
7 3 0 3 1 2 0 3
2 3 3
10 3 0 3 0 1 0 0 1 1 0
2 3 3
11 3 0 3 1 2 2 0 3 0 2 0
4 3 0 3 2
19 3 1 1 0 3 3 0 1 2 3 0 3 1 2 1 0 1 3 0
1 3
18 3 1 1 3 0 2 0 3 1 2 1 1 2 0 3 0 0 3
7 3 2 2 0 1 1 1
11 3 3 2 3 2 1 1 2 0 3 0
5 3 0 3 0 3
3 3 0 3
2 3 3
5 3 0 2 3 0
4 3 0 3 3
3 3 3 0
2 3 1
8 3 0 3 0 3 1 1 0
11 3 3 0 1 2 3 0 0 1 3 0
9 3 3 1 3 3 0 2 3 0
2 3 3
4 3 0 3 0
7 3 0 1 2 2 0 3
2 3 3
5 3 0 3 0 2
7 3 0 3 0 1 2 0
11 3 0 3 1 0 1 2 0 1 1 3
29 3 0 3 0 3 0 3 1 3 0 3 0 3 1 3 1 3 0 0 0 0 1 3 1 0 3 3 3 3
4 3 0 2 3
5 3 0 2 3 0
7 3 3 0 2 2 0 3
4 3 3 1 3
5 3 3 2 0 0
13 3 3 0 1 2 0 3 3 1 3 3 1 3
1 3
8 3 3 0 2 2 1 1 3
20 3 0 3 0 2 1 1 0 1 3 3 2 0 3 3 1 3 1 1 1
2 3 3
10 3 3 0 0 3 3 0 2 1 0
7 3 3 1 1 3 3 0
9 3 3 1 1 0 1 3 3 3
2 3 3
3 3 0 3
2 3 3
5 3 0 2 3 3
3 3 0 3
6 3 3 0 0 1 3
4 3 0 2 3
7 3 1 1 3 3 3 2
3 3 3 3
16 3 3 0 1 1 1 0 2 1 3 3 0 1 3 3 3
2 3 3
7 3 0 3 1 3 3 2
4 3 1 1 3
5 3 3 0 1 0
15 3 3 1 3 2 3 3 3 3 0 3 1 0 1 3
1 3
1 3
5 3 1 1 3 3
5 3 0 2 3 1
7 3 0 2 1 1 3 3
11 3 0 3 3 1 1 1 1 1 3 0
3 3 1 3
4 3 3 0 2
24 3 0 3 0 0 3 0 0 1 3 3 0 1 2 2 0 3 0 2 1 1 2 0 3
3 3 0 3
7 3 0 3 1 3 0 3
4 3 0 3 0
2 3 3
7 3 0 1 3 3 3 0
4 3 0 3 0
3 3 0 3
4 3 2 2 0
19 3 0 3 0 1 3 3 3 1 3 3 1 2 1 1 2 0 3 0
20 3 1 3 1 3 3 0 0 1 3 3 3 0 1 2 1 3 0 0 3
3 3 1 1
12 3 0 1 2 0 2 0 0 1 3 3 0
8 3 0 3 1 3 1 3 0
2 3 3
2 3 3
25 3 3 0 3 3 0 3 1 3 1 3 0 0 1 3 1 3 3 1 3 0 2 0 3 0
2 3 3
2 3 3
8 3 3 1 3 3 2 0 3
16 3 0 3 0 1 2 0 2 3 2 0 1 1 1 2 0
2 3 1
9 3 0 3 1 0 2 0 0 0
16 3 3 1 3 3 3 1 3 3 0 3 0 1 0 2 3
7 3 3 0 1 2 1 3
2 3 3
4 3 0 3 3
7 3 0 3 1 2 2 3
8 3 3 0 2 3 2 0 3
18 3 3 0 1 1 3 1 3 3 3 0 3 3 0 0 1 1 3
7 3 0 2 1 3 0 0
9 3 0 3 1 3 0 0 0 1
4 3 3 3 0
7 3 3 1 3 3 3 0
9 3 0 3 0 3 1 2 3 0
3 3 0 3
4 3 0 3 0
3 3 3 0
11 3 3 0 2 0 3 0 3 3 2 3
7 3 0 3 0 2 1 0
4 3 0 3 2
3 3 1 3
27 3 1 3 1 3 1 3 3 1 2 2 1 3 1 3 3 0 3 0 0 3 0 3 1 3 2 3
9 3 0 3 3 3 0 3 3 2
2 3 0
2 3 3
20 3 0 3 0 1 2 2 0 0 3 1 2 2 0 1 3 3 1 2 0
7 3 3 2 1 0 0 2
3 3 1 3
16 3 0 3 0 2 3 1 2 3 0 0 0 1 2 0 3
4 3 0 3 3
7 3 0 3 0 2 0 3
17 3 2 0 3 1 3 3 0 2 3 0 0 1 3 0 0 0
4 3 0 2 3
2 3 3
6 3 0 3 0 1 2
2 3 3
3 3 1 3
15 3 0 3 1 2 1 2 3 0 1 3 3 3 3 0
20 3 3 1 1 1 1 1 1 1 3 3 3 0 1 1 3 0 0 1 3
3 3 3 0
3 3 0 3
14 3 0 3 1 2 0 3 0 0 1 3 1 3 3
13 3 3 0 0 0 3 3 3 0 1 3 3 1
4 3 1 3 0
4 3 3 0 0
4 3 0 3 3
3 3 1 2
4 3 1 3 0
3 3 3 2
7 3 0 3 0 3 1 0
10 3 3 2 0 0 1 3 0 0 0
3 3 0 1
2 3 3
3 3 0 3
4 3 0 3 3
2 3 3
5 3 0 3 0 0
12 3 0 3 1 2 0 1 3 0 2 0 3
2 3 3
19 3 0 3 0 1 1 3 0 3 0 1 3 3 0 3 0 0 3 0
14 3 0 2 3 1 1 1 2 0 3 1 0 1 2
4 3 3 0 0
2 3 3
7 3 3 1 2 1 3 3
3 3 3 0
4 3 0 3 3
3 3 0 3
3 3 1 3
10 3 3 0 1 1 2 3 1 3 3
4 3 3 0 1
12 3 1 1 1 1 3 0 2 2 0 3 0
2 3 0
4 3 2 0 3
17 3 3 0 1 0 1 2 3 1 0 0 1 3 3 3 3 0
3 3 0 3
13 3 3 1 3 3 3 0 3 3 0 3 0 1
7 3 0 3 1 3 0 3
15 3 0 3 1 0 1 3 3 1 1 1 3 1 1 3
15 3 0 3 1 3 1 0 3 3 3 3 3 0 3 3
6 3 0 3 1 2 3
15 3 3 1 3 3 3 1 3 3 0 1 2 3 1 0
2 3 3
4 3 0 3 0
6 3 0 2 3 0 2
4 3 3 0 0
5 3 1 2 1 3
7 3 1 1 1 1 3 0
3 3 1 0
9 3 3 0 0 3 3 3 0 0
17 3 3 0 0 0 3 3 3 1 0 1 3 2 1 2 0 3
2 3 3
15 3 1 2 0 2 0 1 3 3 0 1 1 3 0 3
9 3 0 3 0 1 0 0 2 3
10 3 3 0 2 2 0 3 0 1 1
1 3
5 3 1 1 3 0
3 3 0 3
2 3 3
4 3 0 0 0
18 3 2 2 3 2 0 3 3 1 2 0 3 0 2 1 3 3 3
3 3 0 2
1 3
6 3 3 0 0 0 1
2 3 3
6 3 0 2 1 3 0
1 3
4 3 3 0 2
3 3 3 0
10 3 1 3 0 0 3 3 3 0 0
2 3 3
4 3 0 3 3
11 3 0 2 1 3 0 1 2 0 3 0
32 3 0 3 0 0 3 1 0 1 3 3 1 2 1 0 1 1 0 1 3 0 0 0 3 3 3 3 1 3 3 0 3
9 3 0 3 1 2 2 0 2 3
11 3 0 3 0 1 2 1 1 2 0 1
4 3 0 3 2
2 3 3
6 3 2 0 1 3 0
7 3 0 3 0 3 0 2
2 3 3
3 3 3 3
6 3 0 3 0 2 0
3 3 0 3
4 3 1 1 1
4 3 0 2 3
1 3
3 3 0 3
2 3 3
3 3 0 3
5 3 3 1 3 0
4 3 0 3 3
31 3 0 0 2 3 0 2 0 3 0 0 1 2 3 0 1 2 0 3 3 0 2 2 2 0 1 0 2 2 2 3
3 3 3 0
14 3 1 3 0 2 3 1 3 3 0 1 1 2 0
3 3 0 3
5 3 0 3 0 2
13 3 1 3 0 2 0 1 3 3 0 3 0 1
3 3 3 2
19 3 0 3 1 2 0 3 0 1 2 0 3 0 1 0 0 1 1 0
11 3 1 1 3 3 0 0 0 0 2 3
6 3 3 3 0 0 0
3 3 0 3
8 3 1 3 0 2 2 0 3
14 3 0 3 0 1 3 3 0 3 1 0 1 3 3
2 3 3
28 3 0 3 0 0 3 1 2 2 3 1 3 1 3 1 3 3 3 1 0 3 1 3 3 3 0 3 3
9 3 1 3 0 0 3 3 0 3
5 3 0 3 1 3
3 3 3 0
8 3 3 1 3 3 3 0 0
4 3 0 3 1
3 3 3 2
2 3 3
3 3 0 3
8 3 0 1 2 1 1 2 3
3 3 3 0
3 3 0 3
2 3 3
4 3 3 0 0
10 3 0 3 1 2 3 0 0 3 3
3 3 3 0
4 3 0 3 3
13 3 0 3 0 3 1 2 1 2 3 1 0 3
25 3 1 3 0 3 3 3 1 2 3 1 3 1 3 0 1 2 3 0 2 1 2 1 3 0
2 3 3
4 3 0 3 0
2 3 3
3 3 3 2
17 3 0 3 3 1 3 3 0 1 3 3 0 3 1 3 1 3
18 3 3 2 0 0 0 1 0 0 3 3 3 0 3 1 2 1 0
3 3 2 3
15 3 1 3 0 0 3 3 1 2 0 3 0 2 0 3
5 3 1 1 1 1
10 3 0 3 0 0 1 3 3 3 0
2 3 3
3 3 0 3
5 3 0 3 1 3
9 3 3 0 2 0 3 0 3 0
4 3 3 2 0
7 3 3 0 2 2 0 3
19 3 0 3 0 1 3 3 3 1 1 1 3 3 0 3 1 1 3 0
5 3 2 0 3 0
22 3 0 3 0 1 1 3 0 3 1 1 3 1 0 3 3 0 1 3 3 1 3
5 3 3 1 2 0
10 3 3 1 3 3 1 2 0 3 0
2 3 3
7 3 0 3 0 3 1 3
8 3 3 1 1 3 2 0 3
3 3 0 2
8 3 0 3 1 2 0 3 0
3 3 3 1
8 3 1 3 0 2 1 1 0
2 3 3
10 3 3 0 1 0 3 3 0 1 2
10 3 3 0 0 0 3 3 3 1 3
6 3 0 2 3 0 0
3 3 1 3
6 3 0 2 3 0 2
2 3 3
4 3 3 0 0
2 3 3
5 3 0 2 3 0
5 3 0 2 3 0
6 3 0 1 0 1 3
3 3 1 1
18 3 3 1 3 3 3 1 3 3 3 0 3 3 0 1 2 1 3
7 3 0 3 0 3 1 3
2 3 3
5 3 3 3 2 0
18 3 0 1 2 1 2 1 3 0 2 0 1 3 3 0 3 1 3
3 3 0 3
22 3 3 1 3 1 1 1 2 1 1 3 1 3 3 0 2 3 0 2 0 2 3
8 3 0 2 3 0 0 1 3
9 3 1 3 0 2 0 2 3 0
8 3 0 3 1 0 1 2 3
3 3 0 3
4 3 2 0 3
15 3 0 3 1 1 1 3 0 2 0 2 0 1 3 3
7 3 0 3 3 1 0 0
2 3 0
2 3 3
9 3 1 1 3 3 3 1 1 3
3 3 0 3
7 3 0 3 1 2 0 3
15 3 0 1 3 3 0 3 1 2 1 1 1 1 3 1
11 3 0 3 0 3 1 0 1 3 3 3
7 3 0 3 0 3 1 2
2 3 3
22 3 0 3 1 3 1 3 1 1 2 0 3 1 2 2 3 1 3 3 0 3 3
5 3 3 1 0 3
3 3 3 2
3 3 3 0
1 3
7 3 0 3 0 3 3 0
2 3 1
21 3 3 0 1 1 1 0 1 3 0 0 3 1 2 2 0 3 1 0 2 0
13 3 0 3 1 2 2 0 3 0 2 0 3 0
6 3 1 1 3 1 2
6 3 0 3 0 2 0
2 3 3
4 3 0 2 3
8 3 0 3 0 2 1 3 0
17 3 0 3 0 2 0 3 1 3 3 1 2 1 3 2 3 3
4 3 0 2 0
10 3 3 1 3 3 3 2 0 0 2
5 3 1 0 0 0
3 3 3 3
3 3 0 3
7 3 1 2 0 1 1 3
17 3 1 3 0 2 0 3 0 0 3 1 2 2 0 2 3 0
2 3 3
8 3 3 0 0 1 2 1 3
1 3
2 3 0
7 3 2 0 3 0 1 1
1 3
6 3 0 0 2 3 0
5 3 3 1 3 3
3 3 1 1
2 3 3
14 3 1 1 1 1 1 3 3 3 0 1 3 3 0
15 3 3 0 2 0 1 3 3 0 3 0 3 3 0 0
1 3
1 3
3 3 0 2
6 3 3 1 3 1 3
2 3 3
2 3 3
2 3 3
10 3 3 0 1 1 1 0 2 3 1
14 3 1 2 0 2 0 1 3 3 3 3 3 0 1
14 3 3 3 0 1 0 1 3 3 3 0 0 1 3
3 3 0 3
5 3 3 0 1 1
4 3 1 3 0
4 3 0 3 3
4 3 0 2 3
7 3 0 3 1 2 0 3
3 3 3 3
10 3 3 1 3 3 0 2 1 0 3
2 3 3
16 3 0 1 3 3 3 1 3 1 0 3 0 0 0 3 3
5 3 2 0 3 0
21 3 3 0 1 1 0 1 3 3 3 1 2 2 3 2 0 1 1 0 0 1
4 3 3 2 0
5 3 0 3 0 3
19 3 3 3 0 2 2 0 3 1 1 1 3 3 1 3 0 2 1 3
3 3 3 2
16 3 3 3 1 3 0 1 1 1 2 3 2 3 2 0 3
7 3 3 0 0 3 0 0
1 3
5 3 1 1 1 1
5 3 0 3 3 0
3 3 3 0
2 3 3
8 3 0 3 0 1 3 3 3
25 3 0 2 1 3 1 2 3 1 3 1 3 3 2 2 0 3 3 1 3 3 0 2 0 3
3 3 1 3
11 3 1 0 1 2 3 2 0 1 2 3
15 3 3 2 1 3 3 3 1 3 3 0 3 1 3 1
15 3 3 2 1 1 1 3 0 0 0 1 2 1 1 3
3 3 3 0
5 3 2 0 0 3
2 3 3
5 3 0 3 0 2
6 3 3 0 0 1 3
13 3 1 3 3 1 2 2 0 3 3 0 1 3
5 3 3 0 1 3
4 3 0 2 3
3 3 3 0
20 3 3 1 1 3 2 0 3 0 2 1 0 3 3 1 0 1 3 3 0
6 3 3 1 0 1 2
6 3 3 1 3 2 0
4 3 0 2 3
3 3 3 2
7 3 0 3 1 3 0 3
11 3 0 3 1 2 0 1 2 0 3 0
6 3 0 2 3 0 1
4 3 1 3 0
6 3 3 0 1 1 1
11 3 3 0 0 0 1 1 3 0 3 0
15 3 3 0 3 3 0 2 3 0 2 3 2 0 0 2
7 3 1 3 1 1 1 1
8 3 0 1 2 1 2 1 2
5 3 0 2 1 3
5 3 0 3 1 3
6 3 3 1 3 3 3
3 3 3 3
11 3 2 0 3 1 3 3 1 1 1 3
8 3 1 1 0 3 3 0 1
3 3 0 3
5 3 0 3 3 0
4 3 0 3 0
9 3 0 3 3 1 3 2 0 0
2 3 0
3 3 0 3
8 3 0 3 0 1 1 0 0
3 3 1 3
5 3 2 0 3 1
2 3 3
4 3 0 3 3
1 3
13 3 1 3 1 3 3 0 3 0 3 0 2 1
12 3 1 3 1 3 3 3 2 0 0 3 3
2 3 3
11 3 0 3 0 1 2 1 3 3 0 0
15 3 0 3 2 0 1 1 3 0 1 1 1 1 1 0
8 3 0 1 0 0 1 0 3
7 3 0 1 1 2 1 3
3 3 1 3
1 3
3 3 3 0
3 3 0 3
6 3 3 1 3 3 3
24 3 3 0 1 2 0 3 1 2 1 2 2 3 0 0 0 3 3 3 0 3 1 3 2
6 3 3 0 1 2 3
6 3 0 1 2 0 2
3 3 1 3
18 3 0 3 3 2 3 3 0 1 3 2 1 1 2 0 2 3 0
16 3 1 3 0 1 1 1 1 2 3 1 3 1 3 1 3
10 3 0 3 1 0 3 3 0 3 0
8 3 0 3 1 3 1 3 3
2 3 3
1 3
1 3
2 3 2
10 3 0 3 3 0 2 0 3 0 3
33 3 3 0 0 1 3 1 3 3 0 3 0 1 1 3 1 3 3 0 0 0 1 3 3 3 1 3 1 3 1 3 0 2
2 3 3
4 3 0 3 0
2 3 3
3 3 3 3
3 3 0 3
12 3 0 3 3 3 0 0 0 0 2 1 3
8 3 3 1 3 0 0 1 3
23 3 0 3 0 3 0 0 1 2 2 0 3 1 3 2 0 1 3 0 2 1 1 3
9 3 0 3 3 1 0 1 2 3
4 3 0 3 3
4 3 3 2 2
4 3 3 0 2
8 3 1 2 0 1 2 0 3
7 3 3 2 0 1 1 3
17 3 1 3 1 3 0 2 0 3 0 1 3 3 0 1 0 3
2 3 3
13 3 0 3 3 1 3 0 1 2 2 0 2 3
11 3 0 3 3 1 3 3 1 2 0 0
2 3 0
3 3 0 3
12 3 0 3 0 1 1 1 1 1 1 0 1
16 3 3 2 0 1 3 3 0 3 1 0 2 0 3 1 3
7 3 0 3 3 0 1 0
16 3 0 2 1 3 0 2 1 1 3 0 1 2 3 3 0
9 3 0 3 1 3 3 2 3 2
14 3 3 1 2 1 2 0 3 1 3 0 1 1 1
3 3 1 0
8 3 1 0 0 1 0 3 3
12 3 0 3 0 2 0 1 2 0 0 3 0
6 3 0 3 0 3 0
2 3 3
10 3 0 1 2 3 0 2 3 0 2
10 3 0 2 3 3 1 3 3 3 3
8 3 1 1 2 3 1 3 1
8 3 3 0 1 1 3 1 3
2 3 3
11 3 0 3 3 3 1 3 3 1 3 0
24 3 0 1 2 2 0 3 1 2 3 0 1 3 2 1 1 1 2 3 1 3 3 1 1
8 3 0 3 1 3 3 0 0
7 3 0 3 2 0 1 3
39 3 0 3 0 0 3 0 0 1 3 3 0 2 3 0 2 0 3 1 2 1 1 2 0 3 1 3 1 3 1 3 3 1 2 0 3 0 0 0
24 3 0 3 0 1 3 3 0 3 0 1 1 0 0 3 0 3 1 0 2 3 1 2 0
3 3 3 3
4 3 3 0 2
4 3 0 3 0
2 3 1
4 3 0 3 3
2 3 3
9 3 3 0 1 1 1 1 1 1
3 3 0 2
3 3 1 3
3 3 3 0
11 3 0 2 3 0 0 0 1 3 0 2
7 3 3 0 1 3 2 1
8 3 0 3 1 2 0 3 0
1 3
3 3 1 3
2 3 3
3 3 3 3
5 3 0 2 3 0
5 3 0 3 1 2
21 3 3 2 0 1 1 2 0 3 0 3 1 2 1 1 2 0 3 0 1 1
2 3 2
2 3 3
9 3 3 1 3 3 3 0 0 3
2 3 3
8 3 0 2 3 0 0 1 3
6 3 1 3 1 3 3
4 3 3 3 2
1 3
10 3 3 3 0 2 0 1 0 3 1
4 3 1 1 3
2 3 2
10 3 0 3 1 3 0 2 1 3 0
9 3 1 0 3 3 3 0 1 0
11 3 0 3 0 2 3 0 0 1 3 0
3 3 3 0
9 3 3 0 0 1 3 3 2 1
9 3 3 1 3 1 3 1 3 3
6 3 3 0 0 1 3
6 3 0 3 0 3 0
28 3 0 2 3 1 3 3 1 3 0 2 3 1 3 3 3 1 3 3 0 3 1 3 0 2 1 3 0
7 3 1 2 0 1 0 1
18 3 0 3 0 1 3 3 0 1 3 3 0 1 3 3 3 2 2
1 3
2 3 0
3 3 3 0
1 3
13 3 1 1 3 3 0 3 3 3 0 3 3 3
5 3 2 0 3 1
2 3 0
1 3
3 3 3 2
22 3 0 3 1 2 1 1 1 3 1 1 3 3 1 2 3 0 3 0 1 2 0
35 3 3 0 2 0 3 0 1 0 3 3 3 2 1 3 3 3 1 1 1 1 1 1 1 2 0 1 1 1 1 2 0 2 1 3
5 3 0 3 1 3
14 3 1 1 1 1 1 3 0 2 1 0 3 3 3
12 3 3 2 3 0 1 3 3 3 1 3 3
11 3 0 1 2 3 0 0 3 1 2 3
3 3 3 0
3 3 0 3
10 3 3 2 3 1 0 3 3 0 3
4 3 3 0 0
17 3 1 3 0 2 2 2 3 1 3 1 3 3 0 3 0 3
7 3 3 1 2 3 1 0
6 3 1 1 3 1 3
22 3 3 0 1 0 1 1 0 1 3 3 1 2 1 2 3 1 3 3 3 0 2
7 3 0 3 1 2 1 0
3 3 0 3
4 3 0 2 3
7 3 0 2 1 3 0 2
12 3 3 0 2 0 3 0 1 3 3 3 0
20 3 0 2 1 3 0 1 0 1 3 0 1 3 0 3 0 3 3 3 0
7 3 0 3 1 2 1 1
9 3 3 1 3 3 0 3 2 3
15 3 3 2 3 1 3 3 0 3 0 3 0 1 3 0
2 3 2
5 3 3 1 3 0
18 3 0 3 0 1 3 3 0 1 3 3 1 0 1 3 3 0 3
16 3 0 3 1 2 2 0 3 0 1 2 3 3 1 3 3
13 3 3 2 3 0 3 0 0 2 0 0 1 2
5 3 0 3 3 0
6 3 0 3 0 2 3
2 3 3
5 3 1 3 2 0
7 3 3 1 0 3 1 1
14 3 0 3 1 0 1 3 3 0 3 1 2 0 3
3 3 1 3
8 3 3 1 3 3 0 0 3
4 3 0 2 3
9 3 0 2 3 0 1 1 3 2
10 3 3 0 2 0 3 0 2 3 0
11 3 1 3 0 1 2 3 1 3 3 0
8 3 3 0 2 0 3 0 3
1 3
6 3 0 3 0 3 0
3 3 3 0
14 3 3 2 1 1 0 1 3 3 3 0 0 1 3
13 3 0 3 0 1 2 1 1 3 2 0 3 0
3 3 1 3
5 3 0 3 3 0
15 3 0 3 1 2 1 2 3 2 0 2 1 3 3 3
8 3 0 3 1 0 1 0 0
8 3 3 0 2 1 2 3 3
2 3 0
4 3 1 1 3
3 3 3 2
1 3
3 3 1 2
15 3 3 0 1 2 3 0 1 2 3 0 3 0 3 3
2 3 1
20 3 0 3 0 2 2 2 3 0 2 0 3 0 1 0 1 3 3 0 3
6 3 1 0 3 0 3
1 3
6 3 0 3 0 0 3
6 3 3 1 3 1 0
6 3 3 1 1 1 1
2 3 3
7 3 2 0 3 0 0 0
2 3 3
3 3 1 3
13 3 3 2 2 3 1 3 3 1 3 3 1 3
9 3 0 0 2 1 1 2 0 3
22 3 3 0 2 0 3 1 2 2 0 3 3 3 0 3 0 3 3 1 3 3 0
6 3 0 0 3 2 3
8 3 0 3 1 3 3 2 0
3 3 1 3
5 3 3 1 2 3
8 3 1 1 2 3 0 0 0
2 3 3
2 3 3
2 3 1
13 3 1 3 0 2 0 3 1 3 0 0 1 3
11 3 0 3 0 1 3 3 3 0 2 3
13 3 0 3 0 1 2 2 0 3 1 0 2 2
4 3 1 2 0
18 3 3 0 0 1 3 0 1 2 3 0 0 0 3 3 3 0 3
2 3 3
7 3 0 3 1 0 1 0
2 3 3
3 3 1 3
3 3 3 0
14 3 3 0 0 3 3 0 1 2 0 3 0 2 3
6 3 0 3 1 2 3
2 3 3
2 3 3
2 3 3
11 3 0 3 1 0 2 0 0 0 1 3
8 3 0 3 0 3 1 3 2
3 3 3 0
11 3 0 1 2 3 1 3 3 0 3 0
12 3 3 1 3 3 1 0 1 3 3 0 3
8 3 3 2 2 0 3 0 0
2 3 1
2 3 3
1 3
2 3 0
8 3 0 1 0 1 0 2 3
8 3 0 3 1 3 1 2 0
1 3
10 3 0 3 1 1 1 1 1 1 3
17 3 0 0 0 2 1 1 1 1 0 2 0 3 1 3 1 3
4 3 3 1 2
15 3 1 3 3 1 3 3 0 3 0 2 3 0 0 3
12 3 0 3 0 1 3 3 0 1 3 3 3
10 3 1 2 1 3 3 0 1 3 1
3 3 3 0
11 3 1 3 2 0 0 1 3 3 1 3
4 3 1 1 3
13 3 0 3 1 2 1 1 1 3 1 3 3 3
10 3 0 3 3 3 3 1 3 3 0
7 3 3 1 3 3 2 3
3 3 1 3
4 3 0 3 3
3 3 1 2
4 3 1 1 3
3 3 3 0
9 3 3 0 1 2 3 0 1 0
3 3 0 3
19 3 0 3 0 1 0 0 2 0 1 2 2 3 1 3 3 2 0 3
3 3 0 3
3 3 1 3
10 3 0 3 1 3 2 0 3 0 0
6 3 3 0 1 0 1
2 3 3
1 3
14 3 3 1 3 0 1 1 1 1 3 2 0 3 0
6 3 0 3 0 2 3
9 3 0 3 0 1 3 3 1 0
3 3 1 3
2 3 3
4 3 0 2 3
1 3
2 3 3
2 3 3
3 3 3 0
15 3 3 0 1 2 1 3 1 3 3 1 2 2 0 3
7 3 3 1 3 3 3 0
2 3 3
15 3 3 1 1 3 0 3 0 1 3 3 0 0 1 2
2 3 1
3 3 1 3
24 3 3 0 0 1 1 1 3 1 3 3 0 1 0 0 1 2 1 1 3 0 1 2 3
6 3 0 3 0 1 2
4 3 0 2 1
5 3 3 2 0 0
5 3 1 1 3 0
4 3 0 3 1
21 3 1 1 3 3 1 3 3 3 0 1 2 2 0 3 1 2 1 0 1 1
6 3 3 0 2 0 1
4 3 0 2 3
9 3 0 2 3 1 3 3 1 3
4 3 3 0 2
8 3 0 3 1 2 0 3 0
8 3 0 3 3 0 1 1 0
4 3 1 1 3
16 3 3 0 2 2 3 1 3 2 3 0 1 3 3 1 3
3 3 0 3
4 3 1 3 0
5 3 0 3 0 2
39 3 3 0 3 3 0 0 3 0 1 2 1 1 2 0 3 3 1 3 3 0 3 1 2 2 0 3 1 3 0 0 2 3 0 0 1 3 0 0
18 3 3 0 2 0 3 0 1 2 1 1 2 0 3 0 1 3 3
7 3 1 3 1 0 3 1
5 3 0 3 1 3
7 3 0 3 1 2 1 0
5 3 1 1 3 3
5 3 2 0 3 0
8 3 0 1 2 1 1 3 1
3 3 0 2
3 3 3 0
31 3 0 2 3 0 2 0 3 1 2 0 3 1 3 3 0 3 2 0 3 0 1 1 1 3 3 3 3 1 2 1
27 3 0 3 1 3 3 0 2 0 3 1 2 1 1 1 0 1 1 0 3 0 1 3 3 3 3 2
21 3 0 3 0 1 3 3 1 2 2 0 2 1 3 1 1 1 1 1 3 0
9 3 3 0 2 1 2 0 1 1
3 3 1 3
3 3 0 2
3 3 0 2
11 3 1 1 3 1 1 1 2 3 2 3
9 3 0 3 0 3 0 2 3 0
20 3 3 3 0 2 1 2 0 1 1 1 1 3 2 0 3 0 1 0 0
3 3 3 0
5 3 1 1 3 0
3 3 0 1
4 3 0 2 3
2 3 3
14 3 0 3 0 1 2 0 1 3 0 2 2 0 3
12 3 1 3 1 3 3 2 1 2 0 2 3
3 3 0 2
4 3 3 1 0
9 3 3 1 3 3 0 1 3 0
6 3 0 1 2 0 3
19 3 0 3 1 2 2 0 3 1 2 3 1 1 1 1 1 1 3 0
2 3 3
2 3 3
4 3 1 3 0
7 3 1 1 1 1 1 3
2 3 3
6 3 3 1 3 3 3
7 3 1 1 3 0 2 3
8 3 0 0 2 3 0 0 0
6 3 0 3 0 2 3
13 3 0 3 0 3 1 0 0 1 0 1 3 3
2 3 3
6 3 3 0 1 2 3
2 3 3
4 3 0 3 0
20 3 1 1 3 0 2 0 3 1 0 2 1 0 1 3 3 1 2 0 3
1 3
1 3
6 3 1 3 0 2 0
5 3 0 3 3 2
13 3 0 3 0 3 1 0 1 0 3 0 3 0
7 3 3 0 0 1 3 0
12 3 1 1 3 3 0 3 1 0 2 1 0
3 3 3 0
3 3 3 2
3 3 0 3
1 3
4 3 0 1 0
1 3
4 3 0 3 3
1 3
26 3 1 3 0 0 3 3 0 3 2 0 3 0 1 2 0 1 0 1 3 0 1 1 1 1 0
3 3 3 0
18 3 1 0 3 3 1 3 0 1 0 1 1 1 2 1 1 1 3
8 3 1 3 0 1 3 0 0
5 3 3 1 3 3
11 3 0 3 1 3 0 3 0 2 1 0
3 3 3 0
1 3
2 3 3
7 3 3 0 2 0 2 1
3 3 1 3
21 3 3 0 3 3 1 3 3 1 2 1 1 1 1 1 1 1 1 1 2 3
17 3 0 3 0 1 3 3 0 0 2 3 0 1 3 3 3 3
8 3 0 3 3 0 2 0 3
14 3 1 1 2 3 0 2 2 0 1 3 0 0 0
7 3 3 0 0 1 3 0
4 3 0 3 2
2 3 0
5 3 0 1 2 3
3 3 1 1
5 3 3 2 0 2
3 3 3 1
3 3 3 0
7 3 2 0 3 0 0 3
16 3 3 1 3 3 3 1 0 0 2 0 3 3 0 0 0
3 3 3 3
3 3 3 0
13 3 3 1 2 1 3 0 1 2 3 1 3 0
12 3 3 1 1 3 3 1 2 1 2 0 1
15 3 3 1 2 2 3 3 1 3 3 1 2 1 0 1
1 3
8 3 0 3 1 2 1 3 1
6 3 0 3 0 3 3
9 3 0 3 0 1 3 3 0 2
6 3 3 1 3 3 3
9 3 0 3 0 1 2 2 0 3
10 3 0 3 1 2 1 3 1 3 3
5 3 0 3 1 3
3 3 0 2
5 3 3 3 0 2
8 3 3 0 1 1 3 0 3
2 3 3
5 3 0 3 3 0
15 3 0 3 1 3 3 1 3 3 0 0 1 2 1 3
1 3
22 3 3 0 1 1 0 1 2 1 0 0 1 3 2 0 1 1 2 0 3 3 0
5 3 0 1 2 1
12 3 3 1 3 3 1 3 3 1 3 1 3
2 3 3
15 3 0 3 3 2 3 0 3 0 2 0 1 3 1 2
21 3 0 2 3 1 1 1 3 1 3 1 3 3 1 2 2 1 3 0 0 0
2 3 3
2 3 0
2 3 1
3 3 3 0
24 3 3 2 0 1 2 1 3 0 0 1 3 0 2 1 3 1 3 3 0 3 1 2 3
9 3 3 0 2 2 3 1 2 2
12 3 3 0 2 3 1 3 3 3 0 2 1
6 3 1 1 3 0 2
11 3 0 3 0 3 0 1 2 0 1 3
3 3 1 2
5 3 0 3 0 2
6 3 0 3 0 1 2
14 3 0 1 1 1 2 0 3 0 1 3 3 1 2
4 3 3 1 0
2 3 0
10 3 0 3 0 2 3 2 0 1 3
7 3 3 1 3 0 3 3
2 3 3
2 3 3
3 3 3 0
6 3 3 1 0 0 3
3 3 1 3
4 3 3 0 1
1 3
3 3 3 0
3 3 1 3
6 3 1 3 1 3 0
7 3 0 3 1 2 0 3
3 3 1 3
5 3 3 1 3 3
1 3
14 3 3 0 1 1 1 2 0 3 0 1 3 3 0
12 3 1 0 2 3 3 0 0 0 0 1 3
10 3 0 3 1 0 0 1 3 3 3
12 3 3 0 2 0 3 1 2 0 1 1 3
7 3 3 1 2 3 3 0
3 3 3 0
3 3 0 3
7 3 3 1 3 3 0 3
1 3
3 3 0 3
19 3 3 1 3 3 1 3 0 3 1 2 3 1 3 3 1 3 3 0
17 3 3 0 0 0 1 1 0 0 2 0 0 2 0 1 3 0
2 3 3
26 3 0 0 2 1 3 0 2 0 3 0 1 3 0 1 3 0 1 2 2 0 3 1 0 2 3
15 3 3 1 3 3 3 1 3 3 1 3 3 1 3 3
9 3 2 0 3 0 1 1 1 3
7 3 3 1 3 3 0 3
3 3 3 2
9 3 0 3 0 3 1 3 1 3
8 3 1 3 0 2 3 3 0
17 3 3 1 3 3 0 3 0 3 0 1 2 1 1 1 1 3
22 3 1 3 0 0 1 3 0 2 0 3 1 0 2 1 2 0 3 0 1 0 0
18 3 3 0 2 1 2 1 3 3 0 2 1 3 3 3 3 0 2
4 3 0 2 3
5 3 1 3 0 0
4 3 0 2 3
14 3 1 3 1 3 3 3 0 2 0 3 1 0 2
11 3 3 1 3 3 0 3 1 3 0 0
2 3 3
7 3 1 3 0 1 1 1
8 3 0 3 0 1 3 3 3
5 3 0 3 3 2
2 3 3
3 3 0 3
2 3 3
17 3 3 1 3 3 0 3 1 0 1 3 3 3 1 0 2 3
3 3 0 1
7 3 1 3 0 0 1 3
1 3
8 3 3 0 2 2 0 1 3
28 3 3 3 1 3 3 0 2 3 1 1 1 2 3 2 0 1 1 1 1 2 1 3 0 2 0 1 2
7 3 1 1 1 1 1 1
14 3 2 0 3 1 3 3 1 0 1 3 3 0 3
2 3 3
18 3 3 1 1 3 3 0 2 0 0 2 0 1 3 3 1 2 3
3 3 3 2
6 3 0 1 2 1 1
20 3 3 3 1 1 3 0 2 3 0 1 0 1 3 3 3 1 0 2 0
7 3 3 1 1 1 1 3
4 3 0 2 3
13 3 3 0 1 1 2 3 1 3 2 0 0 2
7 3 1 3 1 3 3 3
42 3 0 3 1 2 1 2 0 3 0 2 3 2 1 2 0 3 1 3 0 3 0 2 3 1 3 3 0 1 2 1 1 2 0 3 0 2 0 3 0 1 0
12 3 3 3 0 3 3 1 1 1 3 0 0
18 3 0 3 0 2 3 1 1 1 1 3 3 0 1 3 3 0 3
14 3 3 1 3 3 0 3 0 3 1 2 2 1 3
11 3 3 1 3 3 0 3 1 3 0 3
6 3 1 3 1 3 0
9 3 3 1 1 3 2 3 3 2
8 3 0 3 0 1 1 2 3
10 3 0 3 1 2 1 3 2 3 0
3 3 0 3
2 3 3
4 3 3 3 2
5 3 0 2 3 0
3 3 0 3
8 3 1 0 3 3 3 2 0
5 3 0 3 0 3
13 3 1 3 0 2 0 3 3 2 3 1 2 1
10 3 0 1 1 0 1 2 1 3 0
6 3 1 1 3 1 3
5 3 3 0 0 0
1 3
1 3
3 3 0 3
4 3 3 3 2
4 3 3 0 0
3 3 3 0
9 3 1 0 3 3 0 3 3 0
1 3
13 3 0 3 0 1 1 3 0 3 0 1 0 3
3 3 1 2
4 3 3 2 3
21 3 0 3 0 3 1 3 0 3 1 3 0 3 1 3 0 0 1 3 0 0
3 3 1 3
1 3
3 3 1 0
6 3 0 0 2 0 3
7 3 3 1 2 3 1 3
10 3 3 0 0 3 3 0 2 2 1
6 3 3 0 2 3 3
2 3 3
1 3
5 3 1 3 2 0
3 3 0 3
19 3 0 3 1 2 1 2 3 0 3 3 0 3 0 2 2 0 3 0
9 3 3 1 3 3 0 2 0 0
1 3
13 3 1 3 0 2 2 3 0 1 3 3 0 3
4 3 1 2 0
6 3 0 3 0 3 3
11 3 0 3 0 1 0 2 1 1 3 2
2 3 3
9 3 0 3 0 1 3 3 0 2
2 3 1
3 3 3 0
14 3 0 3 0 1 3 3 1 3 3 1 3 3 2
4 3 0 3 0
7 3 1 3 0 2 3 2
31 3 0 3 0 1 1 1 3 3 0 1 3 1 0 1 3 0 2 3 1 3 1 2 0 1 2 0 3 0 2 0
2 3 1
1 3
7 3 0 2 3 0 0 3
5 3 0 3 1 3
7 3 1 3 1 3 3 0
6 3 1 3 0 2 3
16 3 3 1 3 3 0 3 1 2 0 3 0 2 0 2 3
14 3 0 1 2 3 1 3 0 1 1 2 3 2 0
6 3 0 3 0 0 3
2 3 3
2 3 3
3 3 0 3
2 3 3
3 3 0 3
21 3 0 3 0 3 0 1 3 3 0 1 0 1 3 0 1 2 3 1 3 3
11 3 1 3 0 2 0 1 3 3 0 3
18 3 0 3 0 1 3 3 1 2 0 2 0 1 0 0 3 3 3
4 3 3 1 0
2 3 3
11 3 3 0 3 3 0 1 0 1 3 1
4 3 1 2 0
6 3 3 2 3 1 3
6 3 0 2 0 2 3
28 3 0 3 3 1 1 1 2 3 2 0 2 3 0 0 0 1 0 1 3 3 0 3 1 3 3 0 2
8 3 1 3 0 1 2 0 3
3 3 3 0
7 3 1 1 1 3 0 0
2 3 3
2 3 0
19 3 0 3 1 0 1 3 3 0 3 0 1 3 2 0 2 0 1 0
8 3 3 1 3 3 1 2 3
5 3 0 3 0 2
3 3 1 3
2 3 3
8 3 1 3 1 3 0 0 0
1 3
5 3 3 0 0 0
3 3 3 0
2 3 0
12 3 3 1 3 3 0 2 0 1 3 3 2
2 3 3
5 3 0 3 1 3
10 3 0 3 3 1 3 3 0 2 3
4 3 1 3 0
21 3 3 0 1 2 0 3 0 3 0 3 1 0 2 3 1 1 1 1 1 3
5 3 0 3 1 3
17 3 0 3 0 1 0 1 3 3 1 3 1 3 3 3 0 2
7 3 0 3 1 2 0 3
6 3 0 1 3 3 2
3 3 3 0
5 3 0 2 3 0
4 3 3 0 2
9 3 0 3 0 3 3 1 3 1
4 3 1 3 0
4 3 3 2 3
12 3 1 3 0 3 3 3 1 1 3 1 3
2 3 3
8 3 0 0 2 1 3 3 3
1 3
5 3 3 1 0 0
5 3 1 1 3 3
5 3 3 2 0 3
3 3 1 2
2 3 3
11 3 0 3 0 2 0 0 2 3 1 3
9 3 0 3 1 2 2 0 3 0
3 3 0 3
1 3
7 3 0 1 0 1 1 3
2 3 3
3 3 0 3
10 3 0 3 1 0 2 0 0 1 3
1 3
4 3 3 0 0
3 3 3 3
22 3 1 1 3 3 0 1 3 3 0 3 1 3 1 1 3 1 3 3 0 3 0
2 3 3
2 3 3
2 3 3
4 3 0 3 2
7 3 0 3 3 2 0 0
24 3 1 3 0 2 0 3 1 2 2 0 2 3 0 2 1 1 3 0 3 0 1 0 3
8 3 0 3 0 1 3 1 0
23 3 0 3 1 0 2 1 1 3 3 0 1 1 1 1 2 0 3 3 0 0 3 2
11 3 0 3 3 2 2 0 3 1 1 1
5 3 1 3 0 2
5 3 0 2 3 0
3 3 3 3
7 3 3 1 3 3 3 0
3 3 1 2
3 3 0 3
18 3 0 3 0 1 3 3 2 0 1 3 1 1 1 2 0 3 0
6 3 3 0 2 0 3
8 3 0 3 1 3 0 3 3
12 3 3 0 0 1 3 1 3 3 1 2 3
3 3 3 0
4 3 2 0 3
11 3 3 1 1 1 1 3 2 1 1 2
7 3 0 3 0 1 1 3
7 3 3 1 3 3 0 3
1 3
1 3
15 3 0 3 1 2 1 0 2 1 2 0 1 1 1 1
4 3 3 0 0
3 3 1 3
6 3 3 0 0 3 0
1 3
1 3
2 3 3
5 3 0 3 0 3
5 3 3 1 0 0
6 3 0 3 0 2 1
15 3 0 3 3 0 1 1 1 2 0 2 2 0 3 0
7 3 0 3 0 1 3 3
2 3 0
3 3 0 3
3 3 3 0
6 3 3 1 3 2 3
6 3 0 1 0 0 1
17 3 3 1 0 3 1 0 1 3 3 1 0 3 3 0 3 0
11 3 1 3 2 0 2 0 3 1 2 0
4 3 1 0 0
2 3 3
25 3 0 3 0 1 3 3 0 1 0 2 3 1 3 1 3 0 0 2 1 1 1 3 3 0
15 3 3 2 2 0 3 0 2 3 0 0 3 0 2 1
11 3 1 3 0 0 3 3 0 1 2 3
5 3 1 1 3 0
5 3 3 1 3 1
11 3 0 3 0 1 1 3 3 3 0 2
10 3 0 3 0 3 0 3 1 3 3
12 3 0 3 2 0 1 3 0 1 1 0 0
8 3 0 3 0 1 2 0 0
5 3 0 3 0 3
3 3 0 3
2 3 3
4 3 1 0 0
16 3 0 3 0 3 0 3 1 2 2 0 3 1 0 2 1
5 3 3 0 3 3
6 3 0 3 1 3 3
1 3
16 3 1 1 2 3 0 3 0 1 3 3 3 3 1 3 3
4 3 0 2 3
6 3 1 3 0 0 3
19 3 3 1 3 3 3 1 3 3 3 3 3 0 1 3 3 2 0 3
10 3 1 3 0 0 1 3 0 0 0
14 3 3 0 1 1 1 1 0 1 3 0 1 0 0
3 3 1 2
1 3
9 3 0 3 0 0 1 1 1 3
2 3 0
3 3 1 2
9 3 1 3 1 1 3 1 3 1
11 3 3 0 0 1 3 3 0 2 0 1
3 3 0 3
7 3 1 1 3 0 1 0
6 3 1 3 0 1 0
11 3 0 3 3 0 0 3 3 1 1 3
5 3 0 3 0 3
8 3 0 0 2 3 1 1 1
21 3 3 1 3 3 1 3 0 3 0 1 3 3 1 0 1 2 1 1 3 1
3 3 0 3
9 3 0 3 1 2 1 0 1 0
9 3 3 1 0 3 2 2 2 3
2 3 3
4 3 0 3 0
9 3 0 3 0 1 2 1 0 1
6 3 0 2 1 1 3
3 3 0 3
3 3 3 3
3 3 0 1
2 3 3
5 3 0 3 1 2
1 3
18 3 0 3 1 0 1 3 3 1 0 1 3 3 3 0 1 2 3
26 3 0 3 1 2 1 2 0 0 2 3 0 1 1 2 0 2 3 0 1 2 3 0 2 3 2
10 3 3 1 0 1 2 0 3 0 3
2 3 0
9 3 0 3 1 3 0 2 3 0
7 3 0 3 0 1 3 3
5 3 0 2 3 0
14 3 1 1 1 2 0 0 3 3 1 1 1 1 3
3 3 1 3
7 3 0 2 1 1 3 0
11 3 3 1 1 0 3 3 3 1 0 0
9 3 1 3 2 0 2 1 2 3
11 3 0 3 3 1 3 3 0 2 0 0
9 3 3 3 2 1 3 3 0 3
10 3 3 0 1 3 2 2 0 3 0
3 3 3 0
4 3 3 1 0
7 3 3 1 2 3 0 3
1 3
26 3 3 0 2 1 3 0 1 2 3 1 2 1 1 1 3 2 2 0 3 1 2 1 2 0 3
1 3
10 3 0 2 3 0 1 1 2 3 2
4 3 0 3 3
7 3 0 3 1 1 2 3
5 3 3 3 0 2
7 3 0 3 1 0 1 2
8 3 3 1 3 3 2 0 3
7 3 0 3 1 0 1 3
1 3
16 3 1 3 0 2 1 3 1 3 1 1 3 3 0 2 3
11 3 0 3 3 1 3 0 1 3 0 2
1 3
44 3 3 1 0 1 3 3 0 1 1 3 0 2 0 3 0 2 2 2 3 0 1 1 1 1 3 1 1 2 3 0 1 2 0 3 0 3 0 2 1 3 3 0 3
12 3 0 3 0 1 3 3 0 3 3 0 0
12 3 0 3 0 1 3 3 0 3 0 2 3
6 3 3 1 3 0 0
4 3 3 1 0
3 3 3 2
2 3 3
11 3 0 1 2 0 3 1 2 1 1 0
3 3 1 3
3 3 1 3
9 3 0 3 0 1 3 3 0 3
2 3 3
2 3 3
2 3 3
18 3 0 3 0 1 2 3 2 0 3 0 1 2 3 1 3 3 3
12 3 1 3 0 1 1 1 3 2 0 3 0
4 3 0 2 3
6 3 1 3 2 0 0
5 3 1 3 0 0
2 3 3
11 3 0 3 0 1 3 3 1 0 3 3
7 3 0 3 0 3 0 1
3 3 3 0
9 3 3 1 3 3 0 1 3 1
1 3
15 3 1 3 0 2 0 3 3 3 1 3 3 1 3 2
16 3 3 1 3 1 2 1 0 3 0 3 1 2 1 3 0
3 3 1 3
8 3 3 1 0 1 3 3 1
9 3 0 3 1 2 1 1 1 3
12 3 0 3 0 1 3 3 0 1 0 2 1
8 3 0 1 2 1 0 1 3
18 3 3 0 2 2 0 1 3 0 0 0 3 3 3 0 2 0 3
3 3 3 0
6 3 0 3 1 1 3
5 3 3 0 2 0
10 3 3 3 1 3 0 1 3 1 0
6 3 3 2 1 3 3
11 3 3 1 3 3 3 1 3 3 1 3
7 3 3 1 1 1 1 1
7 3 1 3 0 1 1 0
5 3 1 3 0 2
8 3 0 3 1 0 2 3 3
6 3 3 0 0 1 3
4 3 3 1 0
11 3 0 3 0 2 3 0 2 1 2 1
16 3 3 0 2 1 1 3 3 0 1 2 0 1 3 0 2
4 3 1 1 3
19 3 3 1 3 3 1 2 1 2 0 3 1 2 0 1 3 0 0 3
7 3 1 1 3 0 3 3
9 3 3 0 2 0 3 0 1 0
5 3 0 2 1 3
18 3 0 1 2 1 1 1 1 1 1 1 1 3 3 2 0 0 3
23 3 0 3 0 2 3 0 0 1 3 0 0 0 1 3 3 0 1 2 2 0 1 3
4 3 0 2 3
2 3 3
4 3 1 1 3
8 3 3 0 0 1 1 3 0
6 3 3 1 3 3 1
2 3 3
7 3 0 3 1 2 0 3
4 3 0 3 0
3 3 1 3
11 3 1 1 3 0 1 2 3 0 1 0
1 3
9 3 0 2 3 0 1 1 1 0
2 3 3
5 3 0 2 1 3
3 3 0 3
4 3 0 2 3
3 3 3 0
1 3
3 3 0 3
2 3 3
2 3 3
3 3 3 0
3 3 3 0
4 3 0 2 3
2 3 0
3 3 0 3
3 3 0 3
13 3 0 3 0 1 3 3 0 3 0 1 3 3
3 3 0 3
7 3 0 1 3 3 1 3
4 3 2 0 3
3 3 0 3
21 3 0 3 1 3 0 3 1 2 2 0 2 3 0 2 1 3 0 2 0 3
4 3 0 3 3
2 3 3
10 3 3 3 2 0 2 1 0 0 0
25 3 3 0 2 0 3 1 0 1 3 3 3 0 2 0 1 3 3 3 0 1 3 2 3 0
3 3 2 2
8 3 3 1 3 3 0 2 3
3 3 3 2
4 3 3 2 0
17 3 1 3 0 2 3 3 0 2 1 2 3 0 0 0 1 1
1 3
12 3 0 3 1 3 3 1 2 1 1 0 3
5 3 3 0 0 0
2 3 3
17 3 1 1 3 3 1 3 0 2 3 1 2 0 2 0 2 3
4 3 1 1 0
14 3 1 3 1 3 3 0 2 3 1 3 3 0 2
5 3 0 3 3 0
17 3 0 3 0 3 1 0 1 3 3 1 1 3 0 2 3 0
3 3 1 3
4 3 1 1 3
11 3 0 1 3 3 0 1 1 1 1 1
3 3 0 3
2 3 3
5 3 0 3 3 0
4 3 1 3 0
9 3 0 3 0 1 3 3 0 2
17 3 0 2 3 1 3 2 0 1 3 3 3 3 3 0 1 3
3 3 1 3
4 3 0 3 3
3 3 1 3
3 3 3 2
33 3 0 3 0 3 1 3 0 3 1 2 0 0 3 0 2 1 3 2 0 0 1 3 0 2 0 3 2 1 3 3 3 0
14 3 1 2 0 1 2 0 3 1 2 0 0 2 3
2 3 3
10 3 3 0 3 3 0 1 3 1 0
1 3
2 3 3
7 3 2 0 1 3 0 0
5 3 1 3 0 2
19 3 1 2 0 1 3 1 3 3 3 1 2 3 0 2 2 0 3 0
23 3 0 3 1 1 3 1 1 3 0 0 0 1 1 3 3 1 3 0 2 2 0 3
3 3 0 2
10 3 3 0 1 1 1 1 1 0 1
3 3 1 2
18 3 0 3 1 3 1 3 0 2 0 2 0 0 1 3 3 3 3
3 3 1 1
2 3 3
6 3 0 3 0 3 0
15 3 1 3 0 2 2 0 3 1 1 1 3 1 1 3
3 3 1 3
11 3 0 3 0 2 1 1 0 1 2 1
2 3 0
8 3 0 3 0 3 1 2 3
8 3 1 3 3 2 1 2 0
4 3 1 1 3
2 3 3
7 3 0 3 1 2 0 3
8 3 1 0 2 2 1 3 0
9 3 0 3 0 2 0 3 0 2
3 3 1 2
3 3 1 3
13 3 0 3 1 3 3 0 1 1 2 1 3 0
12 3 0 3 0 1 1 3 3 3 1 2 3
9 3 0 3 0 1 3 3 1 3
2 3 3
6 3 3 0 1 1 3
3 3 3 0
3 3 0 3
2 3 3
4 3 1 1 3
2 3 3
30 3 0 3 1 3 0 3 1 2 1 2 0 3 1 2 1 1 3 2 0 3 0 0 0 3 3 3 0 2 0
10 3 0 3 0 3 1 0 1 2 3
17 3 0 3 0 2 0 3 0 2 0 1 2 3 0 1 2 3
14 3 3 1 3 3 0 1 2 3 1 1 1 1 3
12 3 3 1 1 3 3 3 2 3 3 3 0
8 3 0 3 3 0 1 2 3
17 3 0 3 0 3 0 3 3 0 1 3 0 2 0 0 0 3
10 3 0 1 1 1 1 1 1 0 1
3 3 1 3
25 3 0 3 1 2 2 0 3 1 2 1 1 1 1 1 1 1 1 3 3 2 3 0 0 0
8 3 0 3 0 3 1 0 2
6 3 3 2 1 1 2
12 3 0 3 1 0 1 3 3 3 0 1 0
22 3 1 1 3 3 1 3 3 0 2 3 0 0 0 1 0 1 3 3 0 0 3
3 3 1 3
3 3 0 3
9 3 0 3 0 1 3 1 3 3
2 3 3
2 3 3
5 3 0 3 1 3
3 3 1 3
5 3 3 2 1 0
3 3 0 3
15 3 3 1 3 3 1 1 3 3 1 3 3 1 1 3
5 3 0 2 3 1
3 3 3 0
2 3 1
15 3 0 3 1 2 2 0 3 1 1 1 1 1 3 0
6 3 3 1 1 3 3
3 3 1 3
1 3
6 3 0 3 3 1 0
15 3 0 3 0 1 0 2 0 1 1 3 0 1 2 0
2 3 3
2 3 3
13 3 0 2 3 0 0 3 3 1 3 3 2 3
6 3 3 0 1 1 3
5 3 0 3 0 2
6 3 3 0 3 3 3
10 3 1 3 0 1 3 2 0 0 3
6 3 3 0 1 1 3
1 3
3 3 0 3
2 3 3
8 3 3 0 1 2 0 3 0
2 3 3
3 3 0 3
12 3 3 2 0 1 1 2 0 2 3 0 0
3 3 0 3
1 3
7 3 0 3 3 1 3 3
12 3 1 1 3 3 0 3 0 1 0 0 1
7 3 0 3 1 3 0 3
9 3 0 2 3 1 1 1 3 0
7 3 3 0 0 1 2 1
11 3 0 3 0 3 0 1 2 2 0 3
4 3 0 2 3
12 3 2 0 1 3 0 1 0 1 2 1 3
1 3
15 3 3 1 3 3 0 1 3 3 3 2 0 2 0 3
9 3 3 1 0 1 3 3 3 0
15 3 0 3 0 1 2 3 1 3 0 0 3 3 0 3
2 3 3
2 3 3
28 3 3 3 3 2 3 0 1 1 1 1 2 0 3 0 1 3 3 0 1 1 3 0 3 0 2 0 3
2 3 3
3 3 3 0
1 3
4 3 0 3 0
11 3 0 3 0 1 3 3 0 0 3 0
3 3 3 3
6 3 0 1 3 3 3
2 3 3
2 3 3
2 3 0
5 3 3 1 2 3
6 3 3 0 1 1 0
2 3 3
1 3
7 3 0 3 1 0 1 0
3 3 1 3
2 3 3
10 3 3 1 0 1 3 3 0 1 3
6 3 0 3 1 1 3
6 3 0 3 0 1 2
3 3 0 3
3 3 0 3
4 3 0 2 3
4 3 0 3 1
3 3 0 3
1 3
2 3 3
10 3 1 3 3 3 0 2 2 2 3
5 3 1 3 0 2
1 3
4 3 0 3 3
1 3
16 3 0 3 1 1 3 1 3 0 2 3 2 0 3 0 2
3 3 0 3
2 3 3
15 3 0 3 1 2 2 3 2 0 3 0 2 0 2 3
8 3 3 0 2 3 1 3 3
3 3 3 0
12 3 0 3 0 1 2 0 2 2 0 0 3
18 3 0 3 0 1 3 3 0 2 0 0 1 3 3 1 2 1 3
29 3 0 3 1 3 0 2 3 0 2 1 1 1 2 0 0 3 3 1 3 0 3 1 2 3 0 1 0 0
10 3 0 3 0 0 3 3 3 0 3
3 3 3 1
6 3 0 3 2 0 3
3 3 1 3
7 3 3 1 2 0 1 3
3 3 0 3
3 3 0 3
8 3 0 3 0 2 0 0 2
5 3 3 2 0 0
8 3 3 0 1 1 1 0 1
25 3 1 1 3 0 2 1 3 0 2 1 1 3 0 3 0 3 0 3 0 1 3 3 0 3
5 3 0 1 2 3
6 3 0 3 2 0 3
2 3 3
9 3 0 3 0 1 2 1 3 2
9 3 1 3 0 2 1 2 0 3
2 3 3
2 3 3
8 3 3 0 1 1 3 0 0
4 3 3 0 2
3 3 1 3
10 3 3 1 3 3 1 0 1 0 0
26 3 3 1 3 0 2 3 0 1 1 2 0 3 3 1 1 1 3 0 0 3 0 2 0 3 0
3 3 0 3
3 3 0 3
3 3 0 3
5 3 0 2 3 0
3 3 1 3
1 3
5 3 0 3 3 0
8 3 2 0 1 3 1 0 0
13 3 0 3 1 2 3 0 2 1 2 0 2 3
11 3 3 1 2 3 1 3 1 1 0 0
7 3 0 3 1 2 1 1
13 3 0 3 3 1 1 1 1 3 2 2 0 3
2 3 3
7 3 0 1 2 0 1 3
3 3 2 1
6 3 0 3 0 1 2
4 3 0 2 3
2 3 3
9 3 1 1 1 3 1 1 3 0
3 3 3 2
3 3 1 3
12 3 1 1 1 3 2 3 0 2 3 1 3
11 3 0 3 1 2 2 0 3 0 2 3
5 3 3 0 0 3
15 3 0 3 1 2 1 2 3 0 1 3 3 3 0 2
8 3 1 3 0 1 3 2 3
2 3 3
2 3 0
4 3 1 2 3
6 3 0 3 3 2 3
3 3 3 0
12 3 0 3 3 2 3 1 3 3 1 0 2
12 3 0 3 3 0 2 1 1 3 3 0 1
5 3 0 3 0 3
4 3 1 1 1
2 3 3
7 3 3 0 0 2 0 3
6 3 3 2 3 0 3
3 3 0 1
1 3
4 3 3 0 0
8 3 0 3 0 2 0 1 3
7 3 0 3 0 1 2 3
13 3 0 3 1 2 2 0 3 0 1 2 0 3
9 3 3 0 1 1 2 0 2 3
13 3 1 1 3 1 3 0 1 1 1 1 1 0
10 3 1 3 3 0 3 3 3 3 3
4 3 0 3 0
4 3 0 3 0
12 3 0 3 0 3 1 1 3 1 2 0 1
11 3 0 3 1 2 2 3 2 0 2 1
10 3 0 3 0 0 1 0 3 1 1
12 3 1 3 0 2 1 3 0 2 1 1 1
2 3 3
2 3 3
9 3 3 0 2 1 1 3 3 0
4 3 2 0 3
4 3 3 0 0
4 3 0 3 3
8 3 0 3 3 0 2 2 3
12 3 3 1 3 3 0 3 0 1 3 3 2
9 3 1 1 3 0 2 3 2 0
6 3 3 0 1 1 0
3 3 3 0
44 3 3 3 3 1 3 3 1 3 3 0 2 0 0 1 3 3 0 1 3 3 0 3 0 3 0 1 3 3 0 3 2 2 3 0 3 1 3 3 1 3 3 1 3
14 3 3 1 0 1 3 0 2 3 0 1 0 1 3
5 3 0 3 0 3
25 3 3 0 1 1 1 0 2 0 3 0 1 2 1 3 0 1 3 3 0 3 0 1 3 1
3 3 1 2
3 3 0 1
2 3 3
25 3 3 0 3 0 1 3 3 3 1 3 3 0 3 0 3 1 0 1 3 3 0 1 1 3
9 3 3 1 3 0 3 0 0 3
7 3 3 1 1 1 1 0
8 3 0 3 1 3 0 3 0
13 3 0 2 3 0 3 3 3 1 2 1 3 1
21 3 3 1 3 1 0 0 1 3 2 3 0 3 1 2 3 0 0 1 3 0
17 3 1 1 1 3 1 1 2 0 3 0 1 3 3 0 2 3
10 3 3 0 1 1 2 1 2 0 3
8 3 3 1 3 3 1 3 3
9 3 0 3 0 2 3 1 0 3
20 3 3 0 2 2 0 3 0 1 1 2 0 2 3 0 2 0 3 1 3
4 3 1 2 0
3 3 0 1
7 3 0 1 1 3 0 0
3 3 1 3
6 3 3 1 3 3 3
11 3 3 0 2 0 3 1 2 1 1 3
4 3 0 2 3
3 3 1 2
4 3 0 3 3
22 3 0 3 3 0 0 0 1 1 2 1 1 2 0 3 0 3 0 2 3 1 3
5 3 3 3 0 2
10 3 3 1 3 3 0 1 1 3 3
3 3 1 3
2 3 3
11 3 1 1 3 0 2 1 3 0 2 0
1 3
2 3 3
5 3 3 1 2 3
13 3 3 2 0 3 3 0 3 1 1 1 1 1
1 3
1 3
12 3 1 1 1 1 3 2 3 0 1 3 3
6 3 3 1 2 1 3
4 3 2 0 3
1 3
21 3 3 1 3 3 0 3 0 0 3 1 2 1 2 0 3 3 1 2 3 0
2 3 3
16 3 0 2 3 0 1 1 0 1 0 3 0 1 3 0 2
7 3 0 0 2 2 1 3
2 3 3
2 3 3
2 3 3
3 3 1 3
35 3 0 3 3 0 2 2 0 3 0 2 1 3 3 2 0 1 3 0 1 2 3 0 1 2 1 3 0 0 1 3 0 0 1 3
3 3 3 1
2 3 3
38 3 3 1 3 3 3 0 1 2 3 1 3 3 3 1 2 1 2 0 3 3 1 3 3 1 3 0 3 0 0 1 1 3 0 3 0 1 3
10 3 0 3 0 1 2 0 1 3 0
3 3 3 2
6 3 0 3 0 2 3
10 3 3 1 3 3 0 1 3 3 3
10 3 0 3 0 1 0 3 0 0 3
22 3 3 0 1 1 2 0 2 3 0 2 3 3 0 2 0 2 3 1 1 3 3
5 3 3 0 0 0
7 3 3 2 0 1 1 1
8 3 0 1 2 2 0 3 0
4 3 3 0 0
12 3 0 2 3 0 2 0 2 1 3 0 2
4 3 0 3 0
1 3
10 3 0 3 1 1 1 1 1 1 3
2 3 3
2 3 0
11 3 1 0 2 2 3 0 2 1 0 0
10 3 3 1 2 2 1 3 0 0 3
2 3 0
9 3 3 0 2 0 3 0 3 0
6 3 0 1 0 1 3
1 3
11 3 1 3 0 3 3 1 1 1 1 3
3 3 0 3
2 3 3
20 3 0 3 3 0 2 3 1 3 3 2 2 2 1 1 1 2 0 3 3
9 3 0 3 0 2 0 0 0 2
15 3 0 3 3 1 1 1 2 2 0 3 3 0 2 1
4 3 3 1 3
10 3 0 2 3 0 1 1 1 3 3
2 3 3
3 3 3 2
9 3 0 3 0 2 0 3 0 3
4 3 1 1 3
2 3 3
2 3 0
5 3 3 2 0 0
3 3 1 3
5 3 3 1 2 1
3 3 0 3
10 3 3 0 0 2 1 2 0 2 3
9 3 3 0 1 2 0 3 0 2
6 3 0 3 3 0 1
24 3 1 1 3 0 2 0 1 3 3 0 3 1 3 0 0 1 1 3 0 2 2 0 3
7 3 3 0 0 1 1 3
7 3 0 3 3 0 1 3
16 3 1 3 1 3 3 1 3 0 3 0 1 3 1 0 3
3 3 1 3
9 3 0 3 1 1 1 3 1 3
4 3 3 0 2
5 3 0 3 0 2
10 3 0 3 1 1 1 1 3 1 3
7 3 0 3 0 1 3 3
19 3 3 3 1 3 3 3 0 1 1 3 2 1 3 0 0 3 3 1
12 3 1 3 2 0 2 1 3 1 3 0 0
19 3 0 3 0 1 1 1 1 3 1 3 3 3 3 0 0 0 1 0
1 3
3 3 3 0
20 3 0 1 0 1 3 0 2 0 3 0 0 1 1 3 1 3 3 3 2
3 3 3 0
2 3 0
3 3 0 3
5 3 1 3 0 2
2 3 3
8 3 3 1 3 3 0 3 0
19 3 3 1 1 1 1 1 2 0 3 0 2 1 1 0 1 3 3 3
3 3 1 3
1 3
11 3 3 0 2 0 3 0 1 3 3 1
8 3 0 1 0 3 3 1 0
4 3 1 3 0
1 3
15 3 0 3 1 3 1 3 3 3 0 2 0 2 3 0
11 3 0 2 1 1 3 1 3 1 3 0
4 3 3 0 0
3 3 0 1
1 3
11 3 1 3 1 3 0 1 0 1 3 2
3 3 1 0
17 3 0 3 0 1 2 3 3 1 3 3 1 0 1 3 3 3
20 3 0 3 3 0 1 0 2 0 3 0 1 3 3 0 3 0 3 0 1
7 3 0 3 1 3 0 0
2 3 3
5 3 3 1 0 3
3 3 3 2
1 3
3 3 0 3
11 3 1 3 0 1 3 3 3 3 0 3
11 3 3 0 2 3 2 2 2 3 0 1
16 3 3 0 2 0 2 3 0 3 0 1 2 0 3 1 2
1 3
2 3 0
10 3 3 1 3 3 1 3 0 1 3
13 3 3 3 1 3 3 2 1 2 1 1 1 3
2 3 3
2 3 3
11 3 3 0 1 1 1 1 3 0 3 3
6 3 3 0 1 2 3
2 3 3
7 3 0 3 0 1 3 3
8 3 1 2 0 1 2 3 2
5 3 0 3 1 3
6 3 1 3 0 1 3
16 3 2 0 3 0 2 1 3 1 3 3 1 3 1 1 3
4 3 3 0 2
5 3 1 3 0 0
5 3 1 3 0 0
3 3 0 2
8 3 3 1 3 3 0 2 3
23 3 3 1 3 3 3 1 3 3 0 3 0 1 2 0 3 0 2 3 1 0 3 3
28 3 0 1 2 1 3 3 0 1 2 0 1 3 0 2 0 3 0 1 0 1 3 3 1 1 1 1 1
2 3 3
3 3 1 3
11 3 3 0 1 2 1 0 1 2 2 0
14 3 0 3 0 1 3 3 3 0 1 1 0 1 1
3 3 1 3
2 3 3
11 3 0 3 0 1 3 3 0 2 3 0
28 3 3 1 0 1 1 2 0 3 0 1 2 1 2 0 2 3 0 1 1 0 1 3 3 3 1 3 0
3 3 1 3
4 3 3 3 2
5 3 3 1 1 3
10 3 0 3 0 1 3 3 1 3 0
27 3 3 0 1 0 1 3 3 0 3 0 0 3 0 1 3 3 0 2 0 0 1 1 1 2 1 3
2 3 3
15 3 3 2 1 0 2 3 0 3 0 1 1 3 1 1
3 3 0 3
4 3 2 0 3
14 3 1 1 3 0 0 3 0 0 2 0 3 0 3
5 3 1 3 0 1
7 3 3 0 1 1 2 1
3 3 3 3
6 3 3 1 3 0 3
15 3 3 0 2 2 0 3 0 1 0 1 1 2 0 2
5 3 0 3 0 2
6 3 1 3 0 0 0
5 3 3 2 0 0
2 3 3
2 3 3
2 3 3
1 3
9 3 3 1 3 3 0 1 3 3
6 3 3 0 2 0 3
4 3 3 0 0
9 3 3 3 0 2 2 3 0 2
18 3 0 3 0 3 1 3 0 3 0 3 0 1 1 3 3 0 3
1 3
9 3 3 1 2 0 0 1 3 0
9 3 0 3 0 3 1 0 1 2
27 3 3 0 1 0 0 3 3 2 1 0 1 1 1 1 1 1 1 3 1 1 1 1 0 2 0 3
3 3 0 3
3 3 0 3
14 3 0 3 3 0 2 0 3 0 1 3 3 0 3
4 3 3 2 0
8 3 3 1 1 1 1 3 0
2 3 3
8 3 0 3 0 2 1 3 0
6 3 0 3 3 0 2
35 3 0 3 0 1 2 0 1 1 1 1 2 0 3 0 3 0 3 0 1 3 3 0 2 3 3 1 3 0 1 1 1 1 3 1
10 3 1 2 0 3 1 2 1 1 1
4 3 1 3 0
2 3 3
3 3 3 0
13 3 0 3 1 3 0 1 1 2 3 0 0 3
4 3 3 0 2
3 3 0 3
6 3 3 1 3 3 3
19 3 3 0 2 2 0 3 0 2 0 3 1 2 2 0 3 3 1 3
8 3 0 3 0 2 3 0 2
7 3 0 3 1 0 2 0
24 3 0 0 2 3 0 1 1 1 1 2 0 3 0 3 0 2 1 0 0 3 0 3 1
7 3 1 1 3 0 0 0
2 3 0
3 3 1 3
6 3 1 3 0 1 0
2 3 3
1 3
4 3 1 3 2
1 3
3 3 3 0
10 3 1 2 1 3 3 0 3 1 3
2 3 3
18 3 0 3 0 1 0 0 3 2 3 0 3 1 2 1 1 0 1
6 3 1 3 0 0 3
17 3 3 0 2 0 3 1 2 0 3 3 2 2 2 3 0 0
7 3 3 1 2 1 1 1
13 3 0 3 0 1 2 1 2 0 3 1 3 3
3 3 1 0
2 3 0
3 3 0 3
7 3 3 2 1 3 0 0
8 3 0 2 1 3 3 3 3
9 3 0 3 3 1 3 3 3 0
2 3 3
3 3 0 3
3 3 0 3
6 3 1 1 3 0 3
10 3 3 0 0 1 3 0 2 0 3
8 3 3 1 2 2 3 1 2
3 3 3 2
6 3 0 3 0 1 3
3 3 0 1
2 3 3
10 3 3 1 3 3 1 3 0 2 2
5 3 0 3 0 2
3 3 0 3
3 3 3 0
11 3 3 0 1 2 0 1 1 2 1 3
3 3 1 3
1 3
11 3 0 3 0 2 1 3 0 0 1 3
5 3 0 2 0 0
4 3 3 0 0
4 3 0 2 3
4 3 1 3 0
11 3 0 3 1 0 1 0 3 3 3 3
2 3 3
2 3 3
21 3 0 2 3 0 2 0 3 1 2 1 0 2 3 1 3 3 0 1 2 0
1 3
7 3 3 2 0 2 1 2
2 3 3
10 3 1 3 0 1 1 1 1 1 1
12 3 0 3 1 2 1 2 0 1 0 3 0
3 3 3 0
5 3 3 1 0 0
8 3 1 0 1 1 2 1 3
12 3 3 1 3 3 0 2 0 0 0 1 3
5 3 3 1 3 3
6 3 3 2 0 1 1
12 3 0 3 0 1 2 3 0 3 1 1 3
10 3 1 3 0 2 3 1 3 0 0
3 3 3 1
4 3 0 3 0
2 3 0
5 3 1 0 3 3
3 3 3 0
1 3
3 3 1 3
3 3 1 3
17 3 1 3 0 0 3 0 0 2 0 1 2 2 0 3 1 2
3 3 0 3
13 3 3 0 2 1 1 3 1 1 3 3 3 0
12 3 0 3 0 1 2 0 2 3 2 3 0
20 3 0 3 3 1 3 3 0 3 3 3 3 0 1 2 0 3 0 1 2
9 3 3 3 1 3 0 2 0 3
8 3 3 1 3 3 1 0 0
7 3 3 0 1 1 3 3
3 3 0 3
18 3 0 3 1 2 2 0 3 0 2 0 3 0 2 2 0 1 3
1 3
4 3 3 0 0
3 3 1 3
4 3 3 1 3
2 3 3
5 3 0 3 0 3
4 3 1 3 0
4 3 3 0 2
3 3 3 0
3 3 0 1
5 3 1 1 1 2
2 3 3
5 3 2 0 3 0
3 3 0 3
1 3
16 3 1 1 3 3 3 3 3 0 1 3 3 0 1 3 3
3 3 1 2
8 3 0 3 1 3 3 0 0
2 3 3
7 3 0 3 1 3 3 3
2 3 3
22 3 0 3 0 1 3 3 3 0 2 3 3 1 1 1 2 0 2 1 1 3 2
2 3 3
7 3 3 1 3 3 1 2
3 3 1 3
12 3 3 2 0 3 0 1 2 3 1 2 0
3 3 0 3
3 3 1 3
2 3 3
3 3 1 3
16 3 3 0 2 2 0 0 3 0 2 0 3 0 2 1 3
2 3 3
4 3 3 0 0
1 3
7 3 1 3 1 3 3 3
3 3 1 3
5 3 0 3 3 0
7 3 3 0 1 1 1 0
3 3 3 0
19 3 3 2 3 0 1 2 2 0 3 1 2 1 1 1 1 1 1 0
2 3 1
4 3 0 2 3
3 3 1 3
5 3 1 1 1 3
17 3 0 3 0 1 2 0 0 3 3 1 1 3 3 2 1 0
13 3 1 1 3 3 3 0 1 3 3 3 3 3
1 3
1 3
5 3 0 3 1 3
24 3 3 0 2 0 3 0 1 1 1 2 3 1 3 0 1 0 3 3 1 3 1 1 3
13 3 1 1 3 1 3 0 2 0 3 1 2 1
7 3 0 3 0 2 0 3
12 3 0 3 0 1 3 3 3 0 1 1 3
3 3 1 2
2 3 3
2 3 3
16 3 0 3 1 0 1 3 3 0 3 1 3 3 0 2 3
4 3 1 2 3
7 3 0 2 1 3 0 1
6 3 0 3 0 3 0
8 3 3 0 0 1 1 3 0
4 3 1 1 3
6 3 0 3 0 3 3
13 3 0 3 0 1 3 3 0 3 0 2 3 1
6 3 1 3 1 3 0
25 3 0 3 1 2 1 2 3 0 0 0 0 3 3 0 3 0 0 1 1 3 0 2 0 3
7 3 0 3 0 1 0 0
7 3 1 3 1 3 3 0
7 3 0 3 1 0 1 0
6 3 3 1 3 0 3
8 3 3 0 0 1 3 0 0
1 3
6 3 0 3 0 2 3
5 3 3 1 2 3
11 3 3 0 0 1 1 2 0 3 0 1
9 3 3 1 2 1 1 1 1 3
7 3 0 3 0 3 3 0
15 3 0 3 1 2 1 2 0 3 0 3 0 1 2 1
17 3 3 1 3 3 3 1 0 1 2 1 2 0 3 0 3 3
8 3 0 3 1 2 1 1 3
2 3 3
2 3 3
5 3 0 3 1 2
7 3 0 2 1 1 1 3
7 3 3 0 1 2 1 3
6 3 0 3 0 2 3
20 3 0 2 3 0 0 0 1 0 3 0 3 0 1 2 3 1 3 3 3
8 3 1 0 0 3 1 3 0
8 3 0 3 0 3 0 2 3
5 3 3 1 3 3
2 3 3
4 3 3 1 3
17 3 0 3 0 1 2 0 2 0 1 3 0 1 3 3 0 3
2 3 3
5 3 3 1 3 3
1 3
2 3 3
2 3 3
8 3 3 2 1 0 2 0 3
10 3 0 3 0 3 0 1 1 0 1
5 3 0 3 0 3
3 3 3 0
3 3 0 2
5 3 2 0 1 3
1 3
6 3 2 0 3 0 2
21 3 0 3 0 3 0 1 3 3 3 1 3 3 0 3 1 1 1 1 1 2
4 3 0 2 3
9 3 0 3 0 1 2 0 3 0
8 3 0 3 0 1 1 3 3
24 3 0 3 1 3 0 3 0 1 3 3 0 3 3 3 1 3 3 3 1 1 3 3 3
4 3 2 0 3
1 3
1 3
3 3 3 0
2 3 3
5 3 1 3 0 0
4 3 1 0 0
1 3
3 3 1 3
6 3 0 3 0 2 3
31 3 1 3 1 3 3 1 2 3 0 1 2 0 3 0 2 2 3 3 3 1 1 3 1 0 2 3 1 2 0 3
2 3 3
7 3 3 0 2 0 3 0
2 3 3
17 3 0 3 1 3 3 0 2 0 3 0 1 3 3 1 1 3
7 3 3 0 2 0 2 3
3 3 0 3
4 3 3 2 3
1 3
2 3 3
10 3 0 0 3 2 0 3 0 1 3
11 3 0 0 0 1 3 3 3 0 1 0
5 3 3 1 3 3
8 3 3 1 1 3 1 1 3
5 3 0 3 0 2
1 3
5 3 1 3 0 2
3 3 3 1
3 3 3 0
2 3 3
1 3
10 3 1 3 0 1 1 2 0 3 0
5 3 0 3 3 0
4 3 1 2 3
10 3 0 1 2 0 3 1 2 0 3
3 3 1 2
2 3 3
14 3 3 0 1 1 2 0 3 3 1 3 0 2 3
2 3 3
2 3 0
7 3 0 3 1 2 2 0
29 3 1 2 0 2 1 3 1 3 0 3 1 3 1 1 3 3 2 1 3 3 3 3 3 1 3 3 3 3
14 3 0 3 1 2 0 3 3 1 3 3 3 0 0
3 3 3 2
6 3 1 0 0 3 0
13 3 1 0 3 3 0 3 1 2 3 1 3 3
13 3 0 2 3 3 3 3 0 2 3 2 0 3
5 3 0 2 3 0
8 3 3 3 1 3 3 0 2
3 3 0 3
2 3 3
6 3 0 1 2 1 1
12 3 0 3 0 1 3 3 3 1 3 3 3
11 3 0 1 3 3 0 3 0 1 2 3
16 3 3 0 0 1 1 3 1 3 3 3 1 3 3 0 1
3 3 3 0
6 3 3 2 0 0 3
15 3 0 3 1 0 2 0 0 0 1 3 3 3 0 2
6 3 3 1 3 3 3
2 3 3
4 3 3 2 0
3 3 0 3
11 3 1 2 0 2 0 3 1 2 3 1
9 3 0 3 0 2 1 1 2 3
4 3 3 1 0
2 3 3
7 3 0 1 3 3 3 0
1 3
1 3
10 3 0 1 3 3 1 0 2 0 3
15 3 0 3 0 2 0 0 1 0 2 3 1 0 1 3
10 3 1 1 3 3 2 3 1 2 0
1 3
10 3 2 3 1 0 2 2 2 1 3
6 3 0 3 0 1 2
11 3 0 3 1 0 1 3 3 3 0 2
2 3 3
2 3 3
11 3 3 3 1 3 3 3 1 0 1 3
8 3 3 0 0 1 3 3 2
6 3 0 3 1 3 3
2 3 3
3 3 1 3
3 3 0 1
1 3
14 3 1 3 1 3 0 2 3 2 0 1 3 0 2
10 3 0 3 1 3 3 1 3 0 3
12 3 3 0 1 2 3 0 1 1 1 1 3
6 3 3 0 1 1 1
8 3 0 3 0 1 3 3 1
16 3 1 3 0 2 0 1 2 1 1 1 1 1 1 0 2
2 3 3
5 3 0 3 1 3
8 3 0 3 1 2 1 1 0
7 3 0 3 1 3 0 3
7 3 0 1 1 2 3 0
2 3 3
3 3 1 3
2 3 3
3 3 0 3
2 3 3
2 3 2
5 3 3 1 3 3
7 3 0 3 0 1 2 0
4 3 3 1 3
6 3 0 3 0 1 2
19 3 0 3 0 1 3 3 0 3 0 0 3 0 1 2 1 3 0 3
15 3 1 1 3 0 2 0 3 0 1 2 1 1 1 0
3 3 0 3
1 3
2 3 3
19 3 0 3 1 0 1 3 3 1 3 3 3 2 0 2 1 1 3 3
10 3 2 0 3 0 2 1 3 0 0
2 3 3
6 3 3 1 1 1 3
3 3 1 3
2 3 0
8 3 0 3 0 1 3 3 3
6 3 0 3 0 2 0
7 3 0 2 1 3 0 0
14 3 3 0 2 0 1 2 0 1 3 1 3 3 0
7 3 0 3 1 0 2 3
2 3 3
14 3 3 1 3 3 0 1 0 3 3 0 3 0 0
6 3 2 0 1 1 3
10 3 3 1 3 3 1 3 2 0 3
2 3 3
6 3 3 0 1 1 3
1 3
1 3
14 3 1 3 3 0 1 0 0 3 1 3 3 2 0
2 3 3
6 3 1 3 0 2 2
2 3 3
6 3 3 1 3 3 1
3 3 0 3
5 3 0 3 0 3
7 3 0 3 1 2 0 2
17 3 0 2 1 1 2 2 3 1 3 3 0 2 1 3 0 0
27 3 0 2 3 0 2 0 3 1 3 0 3 1 2 1 3 0 2 0 3 3 3 0 3 3 0 3
9 3 3 1 3 1 3 0 1 0
21 3 0 3 0 0 1 3 3 1 2 1 0 2 0 3 0 2 3 2 0 3
2 3 3
8 3 3 1 3 3 1 3 3
10 3 0 3 0 1 3 3 1 3 0
8 3 0 3 0 1 3 3 0
6 3 3 1 3 3 3
2 3 3
2 3 3
3 3 0 3
2 3 3
2 3 3
3 3 3 2
3 3 1 3
16 3 0 3 3 0 1 2 3 2 2 3 1 3 3 1 3
2 3 3
5 3 0 3 0 3
6 3 0 3 1 0 2
4 3 3 3 3
2 3 3
8 3 0 3 0 1 3 3 3
2 3 3
16 3 2 0 3 1 3 3 0 3 0 0 3 1 2 1 0
14 3 0 3 0 3 0 1 3 3 0 2 0 0 3
4 3 1 1 3
14 3 3 1 3 3 3 1 3 3 0 0 3 0 2
2 3 3
12 3 0 3 2 0 3 0 2 0 3 0 0
4 3 0 3 0
4 3 3 0 0
21 3 3 1 3 3 3 0 1 1 1 1 1 0 0 3 1 2 1 1 3 2
9 3 1 3 0 1 2 0 3 3
1 3
13 3 0 2 3 0 1 3 1 3 3 3 1 3
13 3 0 3 3 0 1 2 0 3 3 3 0 1
5 3 3 3 0 2
12 3 0 3 0 3 0 1 3 3 0 1 0
8 3 0 3 0 3 1 2 3
2 3 3
7 3 3 1 2 3 0 0
11 3 0 3 0 1 1 1 1 2 0 3
2 3 3
5 3 0 3 0 3
11 3 0 3 1 0 1 3 3 0 3 0
1 3
14 3 1 1 1 1 0 2 2 1 1 3 0 2 3
22 3 1 1 1 2 0 2 3 1 1 1 2 3 2 0 2 0 3 0 1 3 3
2 3 3
4 3 0 3 0
6 3 0 3 1 3 2
5 3 2 0 3 0
4 3 3 1 2
7 3 3 0 3 1 3 0
7 3 0 3 1 1 1 1
12 3 3 3 1 3 3 0 3 0 1 3 1
10 3 0 3 3 2 1 3 3 1 3
12 3 1 1 3 3 1 2 1 1 1 3 2
6 3 3 1 3 3 0
8 3 0 3 1 3 1 3 3
6 3 0 2 3 0 0
12 3 3 1 3 3 1 0 2 0 0 2 1
21 3 3 2 0 1 0 2 0 1 2 0 1 1 1 1 3 1 3 3 0 3
6 3 3 0 1 1 1
3 3 1 2
3 3 1 3
6 3 0 3 1 2 2
1 3
21 3 0 3 1 0 1 0 1 2 1 3 2 1 2 3 1 1 3 2 1 1
4 3 0 1 2
5 3 1 3 1 3
3 3 0 3
7 3 0 3 0 1 0 3
14 3 0 3 1 2 1 2 3 1 2 1 1 2 3
5 3 3 0 0 0
12 3 0 3 0 1 3 3 0 1 3 3 3
5 3 3 0 1 3
8 3 0 3 1 2 2 0 3
3 3 3 0
2 3 3
29 3 3 2 3 0 3 0 0 3 1 0 1 3 3 1 0 1 1 3 2 1 3 2 3 0 2 0 3 0
4 3 3 0 1
3 3 0 3
7 3 0 3 1 2 0 3
4 3 0 3 0
1 3
9 3 0 3 3 0 2 1 3 3
11 3 3 1 2 1 1 0 1 2 0 0
17 3 3 1 3 0 3 0 1 0 1 3 3 1 2 1 1 3
4 3 0 3 3
13 3 0 3 1 3 0 2 0 2 3 1 0 3
3 3 1 3
3 3 3 0
6 3 3 3 2 0 2
12 3 0 3 1 0 1 3 3 0 3 3 0
3 3 0 1
6 3 0 3 0 3 0
5 3 1 1 0 0
9 3 3 0 2 0 2 3 1 1
12 3 0 2 3 0 1 1 0 1 3 2 1
3 3 3 0
6 3 0 3 0 0 1
4 3 0 2 3
21 3 0 3 0 3 3 0 0 1 2 1 1 2 0 3 0 2 2 0 3 0
5 3 3 0 0 0
7 3 3 0 0 1 3 1
14 3 0 3 0 3 0 1 3 3 2 0 1 3 0
6 3 3 3 1 3 3
2 3 3
2 3 2
4 3 0 2 3
4 3 3 2 0
1 3
3 3 0 3
13 3 0 3 1 2 2 0 2 3 3 1 3 1
9 3 3 1 2 1 1 1 1 1
2 3 3
4 3 3 0 2
2 3 3
3 3 1 2
7 3 1 3 0 0 3 3
5 3 1 1 3 0
2 3 3
11 3 0 2 3 0 2 0 3 3 0 1
12 3 2 0 1 3 0 2 3 2 0 0 2
11 3 0 3 0 1 1 1 3 1 3 0
6 3 0 3 1 2 1
5 3 0 3 1 2
6 3 3 1 3 3 3
1 3
7 3 3 1 3 3 3 0
9 3 0 3 1 2 3 1 2 1
9 3 1 3 1 1 2 0 3 3
7 3 1 1 3 3 1 3
21 3 0 3 0 1 3 3 0 2 3 3 1 3 3 1 2 1 3 0 2 1
2 3 3
13 3 0 3 1 0 1 3 3 1 3 1 3 3
7 3 1 0 3 3 1 3
17 3 0 3 1 2 0 3 0 2 1 0 3 3 0 1 3 3
2 3 3
4 3 0 3 0
11 3 0 3 0 3 0 1 3 3 1 3
2 3 3
3 3 1 3
7 3 0 3 0 0 3 0
7 3 0 3 0 3 1 3
4 3 0 3 0
7 3 3 1 3 2 0 3
9 3 3 3 2 0 2 1 2 3
11 3 1 3 1 3 0 2 3 1 0 3
5 3 0 3 0 3
3 3 3 0
17 3 0 3 3 3 0 0 1 3 3 1 3 0 2 0 2 3
3 3 0 2
2 3 3
6 3 2 3 0 2 3
18 3 3 0 2 1 3 0 0 3 0 3 0 3 3 3 3 1 3
2 3 0
7 3 0 3 0 3 3 0
5 3 3 2 0 0
3 3 3 0
7 3 0 3 0 2 0 3
22 3 3 1 1 3 3 1 2 1 2 0 1 2 1 1 2 1 3 0 2 3 1
29 3 3 3 0 2 0 3 1 2 3 0 1 1 1 2 0 3 1 2 2 0 3 0 1 3 3 0 1 2
4 3 1 1 3
1 3
3 3 0 3
13 3 3 0 1 2 0 3 0 1 3 3 1 2
4 3 1 3 0
5 3 0 3 0 1
3 3 3 0
10 3 0 3 0 1 1 3 1 1 1
1 3
5 3 0 3 0 2
2 3 3
7 3 3 0 1 2 0 3
5 3 1 1 3 0
17 3 3 1 3 3 3 1 3 2 3 1 3 3 1 3 0 2
2 3 3
2 3 0
6 3 1 1 3 1 3
12 3 1 3 0 3 3 3 0 3 1 2 3
12 3 3 0 2 2 0 3 1 3 3 0 3
2 3 3
4 3 1 1 3
8 3 1 1 3 0 3 0 2
2 3 3
12 3 0 3 3 3 1 2 3 1 3 0 0
5 3 3 1 3 3
13 3 0 3 0 1 0 3 3 3 0 2 3 1
3 3 0 3
7 3 0 3 1 2 2 0
13 3 0 3 1 3 3 1 0 2 0 3 0 2
36 3 3 1 3 1 3 0 0 0 1 1 2 1 1 2 0 3 0 1 2 1 3 2 2 3 1 0 3 3 3 3 3 0 1 1 3
4 3 3 0 0
2 3 1
2 3 3
11 3 3 1 3 3 3 1 2 2 0 3
5 3 3 1 3 3
4 3 1 3 0
5 3 0 3 0 3
3 3 0 3
8 3 1 1 2 1 1 0 2
11 3 0 3 0 3 3 3 1 3 1 3
13 3 0 3 1 2 0 0 0 2 0 0 1 2
2 3 3
3 3 0 3
6 3 0 3 1 3 3
15 3 0 2 3 0 1 2 0 3 1 0 1 2 1 0
7 3 2 0 0 3 0 0
7 3 3 2 1 1 3 0
6 3 3 1 0 1 0
4 3 0 3 0
3 3 0 3
2 3 3
5 3 3 0 1 0
4 3 1 3 2
13 3 3 2 1 0 3 1 1 1 0 1 2 3
9 3 3 0 1 1 2 0 2 3
4 3 0 3 0
1 3
13 3 0 3 3 0 1 1 1 1 1 2 0 3
6 3 1 1 3 1 3
1 3
18 3 3 2 0 3 1 0 1 2 1 2 0 3 1 0 1 2 1
2 3 3
8 3 0 1 0 1 1 3 0
2 3 3
5 3 0 3 1 0
1 3
5 3 0 2 3 0
6 3 0 3 0 1 0
2 3 3
25 3 3 1 3 3 0 3 3 0 2 0 3 1 0 2 3 3 2 1 1 3 3 1 3 3
4 3 0 1 0
2 3 3
8 3 3 0 1 1 1 1 0
1 3
11 3 0 3 1 0 2 3 1 0 3 3
26 3 0 1 1 2 3 1 3 3 2 2 0 0 2 0 2 0 0 1 1 2 1 3 2 3 2
3 3 1 3
3 3 3 0
9 3 0 3 0 2 3 3 3 0
9 3 0 1 0 0 2 3 3 0
2 3 3
1 3
4 3 0 3 3
4 3 0 2 3
2 3 3
9 3 0 3 1 2 0 3 0 2
8 3 3 0 2 2 0 3 0
6 3 3 1 0 0 1
4 3 0 1 0
1 3
3 3 3 2
5 3 1 3 0 0
2 3 3
3 3 3 2
15 3 1 3 1 2 3 3 2 0 2 0 3 0 0 3
3 3 3 1
2 3 3
2 3 3
13 3 0 3 1 0 1 0 1 2 2 0 3 0
6 3 0 3 0 1 2
4 3 3 2 1
5 3 0 2 3 0
1 3
9 3 1 1 3 3 0 0 1 3
3 3 3 3
4 3 1 1 3
6 3 3 1 2 3 3
5 3 3 1 3 3
9 3 0 3 1 0 1 3 3 3
4 3 3 0 2
5 3 0 3 3 0
25 3 2 2 0 1 3 3 0 3 0 2 3 0 3 0 2 0 1 3 3 1 3 3 0 3
9 3 3 1 3 3 0 2 3 0
4 3 1 3 0
5 3 0 2 1 3
11 3 0 3 0 1 3 3 1 0 1 3
21 3 0 3 3 1 3 3 3 0 1 2 3 1 3 3 0 3 1 2 3 0
8 3 0 3 0 1 3 3 3
3 3 1 3
3 3 1 3
2 3 3
29 3 0 3 0 1 2 0 1 1 3 0 1 1 2 0 3 0 0 2 1 0 1 3 3 0 2 0 1 3
5 3 3 2 0 3
6 3 2 0 0 1 3
2 3 3
4 3 1 3 0
43 3 3 1 3 3 0 1 1 3 3 3 3 3 3 3 0 1 2 0 3 0 3 0 1 3 3 2 0 1 1 1 0 1 1 0 0 1 0 1 3 1 2 1
1 3
4 3 1 3 0
7 3 0 2 3 1 1 0
13 3 3 1 3 3 0 3 1 0 1 3 1 0
2 3 3
2 3 3
20 3 3 1 3 3 0 1 2 1 1 1 2 0 3 1 3 1 1 3 3
4 3 1 3 0
2 3 3
1 3
2 3 3
6 3 1 3 1 3 1
4 3 3 3 0
3 3 3 0
16 3 3 0 1 2 0 3 0 3 3 1 3 3 1 3 0
9 3 0 0 2 3 1 3 3 3
7 3 0 3 0 3 3 0
3 3 1 3
10 3 0 3 1 2 1 1 2 1 3
26 3 0 3 1 3 3 3 2 0 0 3 3 1 2 2 0 3 0 1 3 3 0 2 1 3 0
4 3 3 3 0
1 3
4 3 3 0 0
1 3
7 3 0 3 3 0 2 2
3 3 3 0
12 3 0 1 0 1 1 1 1 1 3 3 3
2 3 3
7 3 0 2 3 0 1 3
2 3 3
4 3 3 3 0
1 3
3 3 0 3
3 3 1 3
7 3 3 1 3 3 1 3
3 3 1 3
7 3 1 3 2 0 2 0
8 3 0 3 0 0 3 1 2
2 3 0
2 3 3
5 3 0 3 0 2
5 3 0 3 0 2
16 3 0 3 0 1 3 3 3 1 3 3 0 1 3 3 0
3 3 1 1
3 3 1 3
1 3
8 3 3 0 0 1 3 0 2
8 3 1 3 0 2 2 0 3
5 3 1 1 3 3
7 3 3 0 0 1 3 0
20 3 0 3 0 1 0 0 1 1 2 1 1 1 0 1 3 3 3 3 0
2 3 3
3 3 1 3
2 3 3
2 3 3
4 3 0 1 2
37 3 1 1 0 0 1 1 0 2 3 0 1 3 3 0 1 2 0 2 1 2 2 3 0 1 2 1 3 1 3 3 0 1 2 0 3 0
4 3 3 1 0
2 3 3
3 3 1 3
5 3 0 2 3 3
15 3 0 3 0 1 3 3 0 3 0 1 3 3 3 2
1 3
9 3 3 1 3 3 3 1 3 3
19 3 0 3 1 2 1 3 0 0 0 3 3 3 3 1 3 2 3 0
8 3 1 3 0 2 0 1 2
2 3 3
3 3 3 0
11 3 3 0 2 0 1 1 3 0 2 3
1 3
10 3 1 3 0 2 3 1 3 0 3
5 3 0 3 3 0
7 3 0 3 0 1 3 3
4 3 0 1 2
22 3 3 2 0 0 3 0 2 3 0 2 0 3 0 3 0 3 0 2 3 0 2
5 3 0 3 0 3
18 3 0 3 3 0 2 0 2 3 0 2 3 1 3 0 3 0 3
8 3 3 1 0 3 2 1 2
18 3 3 0 1 1 1 1 1 1 1 1 1 2 0 3 0 2 0
2 3 3
11 3 0 3 0 3 0 2 3 1 2 0
4 3 1 3 0
7 3 0 3 1 3 3 3
6 3 3 1 3 3 3
3 3 3 1
31 3 0 3 1 2 3 0 0 3 0 0 2 0 3 0 0 1 3 3 1 2 1 3 2 1 1 1 2 0 3 3
3 3 1 3
10 3 3 0 2 0 3 0 1 2 3
4 3 0 2 3
11 3 3 1 3 3 0 1 3 3 0 3
6 3 0 3 1 3 3
7 3 0 2 0 0 0 0
6 3 0 3 0 2 0
6 3 0 3 0 1 2
4 3 3 0 2
2 3 3
17 3 0 2 1 3 0 2 0 3 1 2 3 0 1 1 1 1
10 3 3 0 0 1 3 1 3 3 0
8 3 3 0 1 2 0 3 0
2 3 3
7 3 1 3 1 3 3 0
20 3 0 0 0 1 3 3 0 3 0 1 3 1 3 3 3 0 0 1 3
7 3 0 2 1 3 3 2
14 3 0 2 2 1 2 2 0 3 0 0 3 0 2
6 3 0 2 3 0 2
3 3 3 0
1 3
1 3
9 3 1 1 3 0 1 1 1 3
12 3 3 1 3 3 0 3 3 1 3 0 0
6 3 1 3 1 3 3
12 3 0 3 0 3 3 2 3 2 0 3 0
8 3 0 3 0 3 1 2 1
1 3
11 3 0 3 3 0 1 0 0 1 1 1
7 3 0 3 0 3 0 1
20 3 0 3 0 3 0 0 1 0 1 3 3 0 1 0 1 3 3 1 1
2 3 3
6 3 0 3 1 3 3
3 3 1 3
10 3 3 2 3 0 1 0 1 1 3
5 3 3 3 0 0
4 3 0 2 3
6 3 3 1 3 0 1
2 3 1
5 3 0 1 2 1
15 3 3 0 2 0 3 0 2 3 3 1 3 3 3 3
6 3 3 1 2 1 3
2 3 1
4 3 3 1 3
7 3 0 3 0 2 3 1
2 3 3
6 3 0 3 3 0 2
11 3 1 2 1 0 3 3 0 3 3 0
12 3 3 0 0 3 3 0 3 1 1 1 2
18 3 3 1 3 3 3 2 3 1 0 3 3 0 1 3 0 2 3
8 3 3 1 3 2 0 3 3
4 3 1 1 3
1 3
17 3 3 0 1 1 1 1 1 1 0 1 3 3 3 0 0 3
23 3 3 0 2 3 1 0 1 3 3 0 3 2 0 3 1 2 2 0 3 3 3 2
4 3 0 3 3
1 3
2 3 3
2 3 3
8 3 0 3 1 2 0 1 3
6 3 0 3 1 3 3
17 3 0 3 1 3 0 3 1 0 1 3 3 1 1 1 3 0
27 3 0 3 0 1 3 3 0 1 3 3 0 3 0 3 3 2 3 2 0 1 3 0 1 2 1 3
23 3 0 3 0 0 3 0 3 1 3 3 3 3 1 3 3 0 1 3 3 0 1 2
13 3 0 3 1 0 1 3 3 0 2 0 0 2
5 3 3 1 3 3
11 3 3 3 1 3 3 3 1 3 0 3
13 3 3 2 0 1 3 0 3 0 1 3 3 3
5 3 0 3 1 3
5 3 0 3 1 2
3 3 1 3
4 3 1 1 1
3 3 0 3
15 3 3 0 0 1 1 3 1 3 3 0 3 1 1 3
1 3
3 3 3 0
6 3 3 0 2 0 3
20 3 3 0 3 3 1 3 1 3 1 1 1 1 1 1 1 1 1 1 1
2 3 3
3 3 0 3
13 3 0 3 0 1 3 3 1 0 1 3 3 3
20 3 3 1 3 3 1 2 1 1 0 0 1 2 1 2 1 1 3 0 1
15 3 0 3 0 1 3 3 1 0 1 3 3 1 2 0
18 3 3 0 1 2 0 3 3 1 3 3 0 3 3 0 2 0 3
3 3 1 2
6 3 3 0 1 1 1
12 3 1 3 1 3 0 1 1 3 2 1 0
3 3 3 0
4 3 0 3 3
5 3 0 3 1 3
4 3 3 2 0
5 3 0 2 3 0
7 3 1 1 3 1 3 3
3 3 1 3
4 3 1 0 3
11 3 0 3 0 3 0 2 3 2 0 3
21 3 1 3 0 2 1 1 1 1 1 3 3 2 3 0 1 3 0 1 1 3
7 3 0 3 1 3 0 3
11 3 3 1 3 3 0 3 0 1 3 3
9 3 0 3 0 1 3 3 3 0
4 3 3 0 2
2 3 3
23 3 0 3 1 2 0 3 0 1 2 0 2 3 1 2 3 0 3 0 1 3 3 3
5 3 0 3 1 3
6 3 0 3 0 3 0
4 3 0 2 3
2 3 3
3 3 0 3
1 3
11 3 3 1 0 1 3 3 1 2 3 0
14 3 0 3 1 3 0 1 1 3 1 3 3 1 2
1 3
6 3 3 0 3 1 0
6 3 1 3 0 1 0
4 3 1 3 0
3 3 0 3
3 3 0 3
5 3 0 3 0 3
4 3 0 3 0
2 3 3
7 3 0 3 1 2 3 0
2 3 3
12 3 0 3 1 0 1 3 3 1 0 2 0
9 3 0 3 3 1 3 3 0 0
5 3 0 3 1 3
18 3 0 3 3 0 2 0 3 0 1 3 3 0 1 1 1 1 3
3 3 3 0
2 3 3
7 3 3 0 2 2 0 3
12 3 0 3 0 1 2 3 0 1 2 3 2
5 3 0 3 3 0
18 3 3 1 3 3 0 3 0 2 0 3 0 0 2 0 2 3 0
2 3 3
7 3 3 0 2 0 2 3
3 3 3 2
7 3 0 3 3 3 3 1
4 3 0 2 3
7 3 3 0 1 1 1 3
14 3 0 2 3 1 0 2 3 1 2 2 0 2 3
8 3 3 0 1 1 1 1 3
11 3 3 0 0 3 3 1 0 1 3 3
6 3 1 3 0 2 1
3 3 0 1
3 3 1 2
4 3 1 3 0
6 3 3 1 3 3 1
5 3 0 3 1 3
4 3 0 2 3
6 3 0 3 1 3 3
3 3 3 0
22 3 3 0 0 3 3 1 0 1 2 1 3 2 0 3 0 1 3 3 3 1 3
2 3 3
3 3 0 3
11 3 0 2 3 1 1 1 3 3 3 3
7 3 0 3 0 2 0 0
6 3 3 0 0 0 1
10 3 0 1 1 3 3 3 1 1 3
10 3 2 0 3 0 2 2 0 3 0
2 3 3
4 3 3 0 2
6 3 3 0 2 3 2
5 3 0 1 2 3
11 3 0 3 1 0 1 2 3 1 2 3
3 3 1 3
9 3 0 3 0 3 3 0 3 3
5 3 0 3 0 3
20 3 3 0 0 0 1 1 0 1 3 3 1 1 3 0 1 1 2 0 1
1 3
3 3 0 3
2 3 3
7 3 3 1 3 3 3 0
2 3 3
5 3 0 3 3 0
19 3 3 1 3 3 3 1 3 2 0 3 1 0 0 1 0 3 0 3
2 3 3
7 3 0 2 3 0 0 0
5 3 0 3 0 1
3 3 0 3
2 3 3
5 3 1 3 0 0
7 3 0 3 3 1 2 2
2 3 3
11 3 1 1 1 1 1 1 3 1 3 0
6 3 3 0 0 1 3
11 3 0 0 3 0 1 0 1 3 3 3
7 3 0 3 1 2 0 2
21 3 0 3 0 3 0 1 3 3 0 3 0 3 0 3 1 3 3 2 0 3
13 3 0 0 0 1 0 1 3 3 1 0 1 3
5 3 1 0 3 3
4 3 3 2 0
8 3 0 3 1 3 0 3 0
6 3 0 3 0 2 1
8 3 0 3 0 0 1 0 0
7 3 0 2 2 1 1 3
16 3 0 3 0 1 3 3 3 1 3 0 3 0 2 3 2
53 3 3 2 0 0 0 3 3 3 1 1 1 1 1 1 1 1 1 3 1 3 0 2 2 3 0 1 1 3 3 3 1 1 0 1 3 0 1 2 3 1 3 1 2 3 3 1 3 3 1 0 1 0
3 3 1 1
9 3 3 0 1 0 1 3 0 3
6 3 3 1 2 1 1
2 3 3
1 3
4 3 1 1 3
12 3 3 1 3 3 0 3 1 2 1 1 0
2 3 3
6 3 3 0 0 1 3
15 3 0 2 3 0 1 1 1 3 2 1 2 3 0 2
5 3 0 3 0 3
30 3 0 3 1 0 2 3 1 2 0 2 3 2 0 2 0 3 0 1 3 3 3 0 0 3 2 3 0 3 0
2 3 0
2 3 3
13 3 0 3 1 2 2 0 3 0 0 0 2 3
10 3 0 3 1 2 1 3 0 2 0
2 3 3
3 3 1 2
2 3 3
1 3
2 3 3
4 3 2 0 3
2 3 1
15 3 1 3 0 1 2 3 3 1 3 3 1 2 0 3
5 3 0 1 0 0
17 3 0 3 0 1 3 3 0 1 1 3 3 3 3 3 2 0
5 3 3 1 0 0
1 3
12 3 1 2 0 2 0 3 1 2 0 1 3
2 3 3
16 3 3 0 0 1 3 1 3 3 0 0 3 1 2 0 3
10 3 0 3 1 2 2 0 3 3 0
8 3 0 3 1 2 2 0 3
11 3 0 3 1 0 2 3 1 3 2 0
6 3 3 0 0 1 3
5 3 0 3 0 2
15 3 1 1 3 1 3 3 3 0 1 2 3 1 3 3
8 3 3 1 3 0 1 3 3
5 3 3 1 3 3
3 3 1 3
3 3 1 3
9 3 3 0 0 1 1 1 3 0
9 3 1 3 1 3 0 0 3 3
1 3
1 3
13 3 3 0 1 3 2 3 0 0 0 0 3 3
12 3 3 2 1 1 3 3 2 0 1 1 3
1 3
2 3 3
4 3 3 1 3
21 3 0 3 0 3 3 3 3 0 0 0 1 3 3 3 0 3 1 0 0 2
4 3 0 2 3
3 3 0 3
13 3 0 3 1 3 1 3 3 0 3 1 2 3
18 3 1 2 0 2 2 3 0 1 2 3 3 0 1 1 2 1 3
18 3 3 1 2 3 0 0 1 3 1 1 1 1 3 1 3 0 2
5 3 3 1 3 3
3 3 3 0
12 3 0 3 1 2 3 1 2 3 1 3 0
10 3 1 3 1 3 3 0 1 0 3
1 3
2 3 3
14 3 0 3 0 1 3 3 1 2 1 3 2 1 0
3 3 1 3
7 3 3 1 3 3 1 2
2 3 3
5 3 3 3 1 2
3 3 0 3
3 3 3 0
1 3
14 3 0 2 3 1 3 3 0 3 0 2 0 0 2
3 3 3 0
9 3 1 2 0 0 3 3 1 3
1 3
18 3 0 3 0 1 3 3 0 3 0 1 2 0 0 1 3 3 2
11 3 1 1 3 1 3 3 0 3 0 3
2 3 3
5 3 0 1 0 0
13 3 0 3 0 1 3 3 3 0 1 2 1 3
12 3 3 0 2 0 3 1 3 0 3 0 2
5 3 3 1 3 3
6 3 0 3 1 3 3
6 3 3 2 1 0 3
3 3 3 0
9 3 0 3 1 2 1 1 1 3
9 3 0 3 1 0 1 0 0 1
3 3 0 3
1 3
3 3 1 3
1 3
5 3 3 1 2 2
5 3 0 3 0 2
4 3 0 3 3
3 3 3 2
3 3 0 3
31 3 3 1 3 3 0 3 1 0 0 3 1 0 0 3 1 0 1 3 1 1 2 0 3 0 1 3 3 0 2 0
4 3 1 1 3
2 3 3
8 3 0 3 0 1 1 1 1
29 3 0 3 0 3 0 3 0 2 0 3 0 1 1 3 3 2 0 3 0 0 0 3 3 2 0 3 3 3
10 3 0 1 3 3 1 0 1 3 3
6 3 0 3 0 2 0
16 3 0 3 0 1 0 3 3 0 3 0 2 0 3 0 1
7 3 2 0 1 3 0 0
4 3 0 2 3
2 3 1
2 3 3
4 3 0 3 3
4 3 3 1 2
5 3 3 0 0 0
3 3 0 3
6 3 0 3 1 0 0
3 3 0 3
18 3 3 1 3 2 2 0 3 0 1 3 3 0 1 2 1 1 3
9 3 3 0 2 0 3 0 3 3
7 3 0 3 1 2 0 3
12 3 3 2 2 2 1 3 0 1 3 2 1
3 3 1 3
1 3
3 3 3 0
2 3 2
5 3 0 3 1 3
10 3 0 1 3 3 1 2 1 0 1
7 3 1 3 0 1 0 3
11 3 3 0 2 0 3 0 1 2 0 3
1 3
3 3 0 1
5 3 1 3 0 0
1 3
6 3 1 1 3 3 0
10 3 0 3 0 3 0 1 3 3 3
11 3 3 0 2 3 2 0 2 2 0 3
13 3 0 2 3 0 3 1 3 3 0 0 2 0
3 3 0 3
5 3 0 3 3 0
3 3 3 0
9 3 3 3 0 0 0 3 3 3
28 3 0 1 0 1 3 3 0 1 2 3 0 1 3 2 1 2 0 3 0 3 1 1 3 3 0 3 0
18 3 1 1 3 1 3 1 3 0 0 1 2 1 2 1 1 1 3
11 3 0 3 0 3 0 1 3 3 1 3
12 3 3 2 0 1 1 2 0 3 1 3 3
8 3 3 1 3 3 3 0 0
2 3 1
5 3 3 2 1 0
2 3 3
2 3 0
17 3 0 3 0 3 0 1 3 3 3 1 1 3 3 0 2 3
3 3 3 2
3 3 1 3
4 3 0 2 0
5 3 3 2 0 2
3 3 3 2
7 3 0 0 2 3 0 0
2 3 3
2 3 3
22 3 0 3 1 0 1 3 3 1 2 1 1 1 3 3 3 3 1 2 0 2 0
4 3 0 2 3
4 3 0 2 3
6 3 0 3 1 3 3
2 3 3
6 3 1 3 1 3 3
1 3
4 3 0 3 0
7 3 1 1 1 3 1 3
3 3 3 0
6 3 0 1 0 1 3
4 3 1 3 0
3 3 3 0
4 3 2 0 3
3 3 1 3
2 3 3
3 3 1 2
3 3 0 3
5 3 0 3 0 1
2 3 2
5 3 0 3 1 2
2 3 1
3 3 0 2
35 3 0 2 1 3 0 2 1 2 2 3 1 3 0 2 3 0 2 0 3 0 3 1 2 3 1 3 3 0 1 0 2 3 3 1
3 3 3 0
4 3 0 1 1
2 3 3
23 3 2 1 0 3 3 3 3 3 0 0 0 1 3 3 1 3 1 3 1 3 3 3
3 3 3 2
3 3 3 2
7 3 0 3 0 2 1 3
2 3 3
3 3 0 3
3 3 0 3
5 3 3 0 1 0
9 3 3 1 3 3 1 3 0 3
4 3 1 0 3
8 3 3 0 0 0 3 0 2
4 3 2 0 3
9 3 1 3 0 2 2 0 3 1
14 3 3 0 1 1 1 0 1 3 3 3 0 3 3
7 3 3 1 3 3 3 0
2 3 3
2 3 0
1 3
5 3 3 0 2 0
3 3 1 3
2 3 3
7 3 0 3 1 2 3 0
9 3 3 1 3 0 2 3 0 0
2 3 1
2 3 3
11 3 0 3 0 1 3 3 3 0 1 0
3 3 3 0
5 3 3 1 3 0
6 3 3 0 2 0 2
3 3 0 3
2 3 3
2 3 1
7 3 3 3 1 3 0 3
2 3 3
9 3 0 3 1 2 2 1 3 0
3 3 0 3
17 3 3 0 1 1 2 3 1 3 3 1 2 2 1 1 3 0
19 3 1 1 3 1 3 3 0 0 1 1 1 0 1 3 3 3 0 3
3 3 3 0
2 3 0
12 3 1 3 0 1 2 3 0 0 0 1 2
7 3 0 3 1 3 3 2
13 3 1 3 0 0 3 3 1 1 1 1 2 0
3 3 3 0
9 3 3 1 3 3 0 3 1 2
2 3 3
3 3 0 3
2 3 3
8 3 3 1 3 3 3 3 0
4 3 0 2 3
3 3 3 0
3 3 0 3
4 3 1 3 0
3 3 1 3
8 3 0 3 0 1 2 3 3
6 3 0 3 0 1 0
8 3 0 3 1 1 3 0 0
6 3 0 3 0 3 3
7 3 0 1 3 3 1 2
2 3 3
13 3 0 3 0 1 3 3 0 1 0 2 1 0
8 3 0 3 0 1 2 0 3
4 3 2 0 3
13 3 0 3 0 1 3 3 3 0 2 1 3 2
7 3 3 1 2 1 0 1
3 3 0 3
3 3 1 3
5 3 0 3 0 3
1 3
4 3 0 3 0
3 3 3 0
9 3 2 3 0 1 2 3 0 2
10 3 2 0 3 0 2 2 0 3 0
9 3 1 3 0 0 1 3 0 0
5 3 2 0 3 0
23 3 0 3 1 2 3 0 0 1 3 0 2 0 1 3 3 3 0 1 2 0 3 3
3 3 0 3
4 3 3 1 3
2 3 3
12 3 0 1 3 3 0 3 0 2 0 1 3
16 3 0 2 3 0 2 0 0 2 0 1 1 3 1 3 0
9 3 0 2 3 0 2 0 3 0
13 3 1 3 0 1 2 0 3 0 1 0 0 2
7 3 3 1 3 3 1 3
11 3 3 0 0 0 1 0 1 2 0 2
4 3 1 3 0
1 3
18 3 1 3 0 2 0 3 0 1 2 0 3 0 2 0 1 3 3
2 3 0
12 3 0 3 0 1 3 1 3 3 0 1 3
4 3 3 0 1
4 3 1 0 0
8 3 3 0 1 2 0 3 0
2 3 3
3 3 3 0
6 3 2 0 3 1 3
5 3 0 3 0 2
1 3
6 3 3 0 0 1 3
5 3 0 3 0 2
1 3
4 3 0 3 3
9 3 3 1 1 1 1 1 1 1
4 3 2 0 3
25 3 0 1 3 3 0 1 3 3 0 3 0 2 2 3 3 3 1 2 1 1 0 1 2 3
23 3 1 3 0 2 0 3 0 3 1 3 3 3 0 3 1 2 1 3 1 3 0 0
1 3
13 3 0 3 0 1 1 1 1 3 3 3 0 3
9 3 3 1 3 3 0 3 0 3
12 3 3 0 1 1 1 1 2 0 3 0 2
4 3 3 3 0
4 3 0 3 3
3 3 0 1
3 3 1 3
6 3 3 0 0 1 3
5 3 0 3 3 0
7 3 3 0 1 1 1 3
15 3 3 0 1 1 0 1 3 3 3 3 1 3 3 3
9 3 1 3 1 3 3 1 3 0
3 3 0 3
12 3 3 0 0 0 3 3 3 0 1 3 0
4 3 0 2 3
13 3 1 3 0 2 3 2 0 0 0 3 3 1
11 3 0 3 3 1 1 1 1 1 3 0
3 3 3 0
7 3 3 0 2 1 2 3
1 3
5 3 0 3 1 3
11 3 0 3 3 1 3 3 0 3 3 3
2 3 3
6 3 0 1 1 2 3
5 3 2 0 3 0
3 3 0 2
2 3 3
17 3 0 3 1 2 1 1 0 1 3 3 3 2 0 1 3 0
3 3 0 3
4 3 0 2 3
4 3 2 0 3
10 3 0 3 3 0 1 1 2 0 3
6 3 3 0 0 1 3
6 3 1 1 3 1 3
15 3 0 3 1 2 1 1 2 0 3 0 1 2 3 3
6 3 3 3 3 0 1
6 3 0 3 0 1 0
3 3 3 0
2 3 3
3 3 3 0
17 3 0 3 1 3 3 0 1 1 2 0 3 0 3 1 1 3
12 3 3 1 3 3 0 1 2 1 1 1 0
2 3 0
4 3 1 3 0
9 3 3 0 2 1 3 1 3 3
9 3 0 3 3 1 1 3 1 3
3 3 3 2
2 3 3
37 3 3 0 1 2 3 0 3 1 1 1 1 1 1 1 1 1 1 1 1 3 1 1 2 0 3 0 3 1 2 3 0 0 1 3 0 2
10 3 1 3 1 3 1 2 0 2 0
16 3 0 3 0 1 1 0 2 3 0 1 3 3 0 3 3
4 3 1 3 0
3 3 1 3
2 3 0
21 3 0 3 3 0 2 0 1 2 3 0 2 0 3 1 2 0 0 0 1 3
5 3 1 1 3 3
9 3 0 3 1 3 0 3 0 3
17 3 3 1 1 0 3 0 2 0 1 2 1 1 1 1 1 0
2 3 3
14 3 3 0 1 1 3 0 1 0 3 0 1 3 3
10 3 0 3 0 3 1 2 1 2 0
2 3 3
2 3 3
7 3 3 1 3 3 3 0
3 3 3 0
4 3 0 1 0
9 3 0 3 1 3 3 1 0 2
1 3
3 3 1 3
30 3 0 3 3 1 1 2 1 3 0 0 3 3 0 1 1 3 0 2 3 0 0 1 3 0 0 1 3 0 2
2 3 3
4 3 3 2 1
2 3 1
22 3 0 3 0 3 1 2 1 1 1 2 0 3 0 1 3 3 0 3 1 2 3
5 3 1 3 0 0
21 3 3 1 3 3 0 2 0 3 1 3 0 3 3 0 0 1 3 0 0 1
7 3 3 1 3 0 2 3
5 3 0 1 0 0
3 3 3 3
24 3 0 3 0 3 1 0 1 3 3 0 0 3 0 0 3 1 2 1 1 2 0 2 0
2 3 0
3 3 0 3
2 3 0
16 3 0 1 2 0 3 0 1 2 3 1 3 0 1 0 1
4 3 1 3 2
6 3 0 3 3 3 3
4 3 3 0 0
3 3 3 2
19 3 2 0 3 0 2 1 3 0 1 1 2 0 3 1 3 3 3 2
4 3 3 3 1
1 3
3 3 1 3
3 3 3 1
1 3
4 3 1 3 0
17 3 3 1 3 3 0 1 0 1 0 1 2 1 2 0 2 3
3 3 3 0
3 3 3 3
2 3 3
2 3 3
6 3 3 0 0 0 1
4 3 1 3 0
6 3 0 3 1 2 3
3 3 3 0
3 3 1 2
10 3 3 0 1 1 2 3 1 3 3
2 3 3
3 3 3 1
25 3 0 3 0 2 1 1 2 1 1 2 3 3 3 3 2 0 2 0 2 1 1 3 0 0
9 3 0 3 0 1 3 3 0 3
2 3 3
8 3 0 3 3 0 2 0 3
13 3 0 1 3 3 3 3 1 0 2 3 0 3
5 3 1 0 3 3
4 3 3 0 0
3 3 3 3
3 3 0 3
2 3 3
3 3 3 0
2 3 3
1 3
6 3 3 0 2 3 2
11 3 0 3 0 1 3 3 0 1 0 3
8 3 0 3 1 2 1 2 3
5 3 3 0 0 0
24 3 3 0 2 0 3 3 1 3 3 1 0 0 2 1 1 3 3 1 3 3 1 1 2
3 3 3 0
3 3 1 3
6 3 0 2 3 0 3
2 3 3
2 3 3
8 3 2 0 3 0 2 0 3
6 3 3 0 2 0 3
1 3
5 3 1 1 3 3
5 3 2 0 1 3
2 3 3
7 3 0 3 1 3 1 3
7 3 3 1 2 0 3 0
4 3 1 1 3
3 3 0 2
13 3 1 1 3 1 3 3 1 2 1 1 1 3
4 3 0 3 3
3 3 3 0
3 3 1 3
2 3 1
5 3 1 3 0 2
10 3 0 3 1 0 1 3 3 0 3
3 3 1 3
22 3 1 3 0 2 1 1 1 3 0 1 0 0 3 1 0 1 3 3 1 0 0
3 3 0 3
7 3 0 0 0 0 2 0
25 3 3 0 0 1 3 0 0 3 3 1 2 0 3 1 3 0 3 0 1 2 2 0 3 0
6 3 2 0 3 0 1
14 3 3 1 1 3 3 3 0 3 1 3 3 0 3
2 3 3
4 3 0 0 1
13 3 1 3 0 2 1 2 0 2 1 3 0 1
2 3 3
4 3 0 0 1
3 3 3 0
10 3 0 3 1 3 0 2 0 3 3
1 3
3 3 3 0
2 3 3
11 3 0 3 1 2 1 2 0 3 0 3
15 3 3 1 3 3 3 0 2 2 0 3 0 0 1 3
2 3 3
3 3 0 3
2 3 3
4 3 2 0 3
2 3 3
24 3 1 3 3 2 2 0 3 0 0 3 0 1 1 1 1 1 3 0 1 1 2 1 0
7 3 3 1 3 3 3 0
13 3 0 3 3 1 2 3 0 2 3 0 1 0
9 3 0 3 1 2 0 3 0 2
9 3 0 3 0 0 0 2 3 0
1 3
4 3 2 0 2
10 3 0 3 0 3 1 2 2 0 2
3 3 0 3
4 3 0 2 3
6 3 3 3 0 0 0
10 3 1 1 1 3 0 1 3 3 3
6 3 1 3 1 3 3
5 3 1 1 1 3
8 3 0 3 3 0 3 3 3
4 3 1 1 3
8 3 0 2 3 0 2 2 2
6 3 3 0 0 1 3
1 3
1 3
44 3 1 0 3 3 1 1 2 2 1 0 1 3 3 0 3 1 0 3 3 0 3 1 2 0 3 0 0 1 3 0 0 0 3 3 3 3 2 0 0 1 0 1 3
2 3 3
8 3 3 0 2 2 0 1 3
11 3 1 3 0 1 1 3 0 1 3 3
3 3 0 3
2 3 2
9 3 3 0 2 1 0 2 1 3
1 3
4 3 3 1 0
18 3 1 3 0 1 1 3 2 3 0 1 3 3 3 3 0 1 3
3 3 3 2
4 3 0 3 0
6 3 0 3 1 3 0
9 3 3 0 1 2 3 1 2 3
1 3
14 3 0 3 0 1 3 3 0 3 1 1 1 1 0
3 3 0 3
4 3 0 3 0
4 3 3 2 0
9 3 1 1 1 1 3 0 3 2
1 3
5 3 3 1 3 3
2 3 3
3 3 1 3
8 3 3 1 3 3 1 3 0
12 3 0 3 1 3 0 2 0 2 3 0 3
4 3 0 2 3
7 3 0 1 1 1 1 0
8 3 3 1 3 3 3 0 3
24 3 0 3 1 1 3 1 3 0 2 1 3 0 0 0 2 2 0 3 0 2 2 0 3
3 3 3 2
11 3 0 3 1 2 1 3 3 1 1 3
3 3 1 3
3 3 0 3
17 3 3 1 3 3 1 1 1 3 0 2 0 3 0 3 0 3
6 3 1 3 0 1 0
9 3 0 3 1 0 1 3 3 3
1 3
2 3 3
19 3 0 3 1 2 0 3 1 1 1 3 2 1 2 0 3 0 2 1
7 3 3 1 3 3 3 1
5 3 1 1 3 0
6 3 3 0 2 3 3
10 3 1 1 1 3 3 0 1 3 3
2 3 3
3 3 3 1
5 3 1 0 0 0
5 3 3 1 3 3
9 3 0 2 3 0 1 1 3 2
4 3 0 2 3
4 3 1 3 0
4 3 0 2 3
5 3 0 0 1 2
8 3 0 3 1 2 3 0 2
4 3 0 2 3
13 3 1 3 0 0 0 1 1 3 0 3 1 3
17 3 3 3 1 1 3 0 1 1 2 3 0 1 3 3 3 0
12 3 3 2 0 2 0 3 3 0 0 3 3
5 3 3 0 2 1
2 3 3
6 3 0 3 0 2 0
12 3 0 3 1 3 0 2 3 0 1 1 0
18 3 0 3 0 1 2 1 1 2 3 1 3 3 1 0 1 3 3
9 3 0 3 0 3 1 2 0 3
6 3 3 0 0 3 3
9 3 3 0 2 0 3 1 3 0
3 3 3 3
29 3 0 3 0 2 2 0 2 2 0 3 0 2 0 3 0 0 3 0 0 3 1 2 1 1 2 0 3 0
17 3 0 3 1 2 1 2 0 3 0 3 0 3 0 2 3 0
17 3 0 3 1 2 1 2 3 2 0 3 3 3 3 2 3 0
21 3 3 1 1 2 1 1 1 1 1 1 1 1 1 3 3 3 2 1 3 0
17 3 3 0 0 1 3 1 3 3 0 3 3 1 0 1 2 3
15 3 0 0 2 0 2 0 1 1 1 1 0 2 0 3
8 3 1 3 0 1 2 1 3
3 3 3 1
6 3 3 0 2 3 3
12 3 0 3 0 2 0 0 2 0 2 1 3
5 3 3 1 3 3
2 3 1
3 3 1 3
7 3 0 3 1 0 2 0
8 3 3 1 3 3 3 1 2
3 3 0 3
30 3 3 1 3 3 3 1 2 0 1 3 1 3 3 1 2 0 3 1 3 3 0 1 3 3 0 2 3 0 3
1 3
6 3 0 3 0 1 0
9 3 1 3 0 0 0 1 1 2
2 3 3
7 3 0 3 3 0 0 0
7 3 3 0 1 2 0 3
3 3 0 1
11 3 0 3 1 0 1 3 3 1 2 3
4 3 0 3 3
1 3
3 3 1 3
7 3 0 3 1 3 1 3
20 3 1 3 0 0 1 3 0 1 2 0 3 0 3 0 3 1 2 1 3
5 3 1 1 3 3
10 3 3 0 3 2 0 0 3 0 0
5 3 0 2 3 0
12 3 0 3 0 1 3 1 1 1 1 1 0
8 3 3 1 3 3 3 0 2
10 3 0 3 0 3 0 3 1 3 1
8 3 3 3 0 2 3 3 0
6 3 0 3 0 2 3
2 3 3
12 3 0 3 0 2 0 0 2 0 3 1 2
9 3 0 3 0 1 3 3 0 3
17 3 0 3 1 2 2 0 3 1 0 2 0 1 2 1 3 0
8 3 1 3 1 0 1 2 3
8 3 3 1 2 0 1 1 3
8 3 3 1 1 1 3 3 3
5 3 3 0 1 3
11 3 0 2 3 0 0 0 1 1 3 0
17 3 0 3 1 3 1 3 3 0 3 1 3 0 1 2 1 3
7 3 0 3 3 1 3 3
3 3 3 0
6 3 0 1 3 3 3
6 3 0 3 0 3 3
12 3 0 3 1 3 3 0 2 0 3 1 2
4 3 0 3 3
7 3 3 0 1 1 1 0
4 3 3 2 3
8 3 0 3 0 1 3 3 3
3 3 0 3
8 3 0 3 1 1 3 1 3
17 3 0 3 0 3 3 1 3 3 3 1 0 2 0 2 3 2
5 3 2 0 3 0
1 3
5 3 0 3 1 0
2 3 3
7 3 3 0 1 1 1 3
3 3 3 3
3 3 0 3
10 3 3 0 1 2 0 3 0 3 2
24 3 3 1 2 0 3 0 2 1 1 3 0 1 3 3 3 3 1 2 3 0 3 0 3
9 3 0 0 2 3 0 1 1 0
1 3
2 3 3
10 3 3 1 3 3 3 1 3 3 3
15 3 0 3 0 1 0 0 1 3 3 3 1 2 0 3
7 3 0 3 3 0 2 0
6 3 0 3 0 2 3
2 3 3
32 3 0 1 1 3 3 3 0 3 0 1 3 3 3 0 3 3 0 1 3 3 0 3 1 0 1 2 2 3 2 3 3
4 3 0 3 0
1 3
2 3 3
5 3 3 1 3 3
3 3 1 3
9 3 0 3 0 0 3 1 2 3
2 3 3
5 3 3 0 0 3
3 3 3 0
15 3 3 1 3 3 0 1 3 3 3 0 0 0 1 0
4 3 1 2 0
25 3 3 2 1 1 2 0 3 0 1 1 2 3 1 2 3 0 3 1 3 1 3 0 0 3
8 3 0 3 1 2 1 1 3
1 3
20 3 0 3 0 1 2 3 3 1 3 3 1 3 0 2 0 3 1 1 3
6 3 3 3 0 3 3
4 3 0 3 3
7 3 0 3 1 2 3 0
3 3 1 3
2 3 3
3 3 3 0
7 3 0 3 1 1 1 3
6 3 0 1 2 3 0
7 3 3 0 0 1 3 0
16 3 0 3 1 3 3 0 1 1 2 3 1 3 3 0 3
5 3 3 0 2 2
3 3 0 3
9 3 0 3 1 3 3 1 2 3
21 3 3 1 3 3 0 1 0 0 1 3 3 3 3 1 3 3 3 1 3 1
2 3 3
3 3 0 3
4 3 0 3 3
11 3 3 0 0 1 3 0 1 2 2 3
3 3 3 2
4 3 0 3 0
22 3 3 0 1 1 1 2 0 3 0 3 1 3 1 1 1 1 3 0 3 3 3
3 3 1 3
8 3 0 2 3 0 2 0 3
18 3 0 1 1 2 0 3 1 1 1 1 1 3 0 0 1 3 0
7 3 0 3 0 3 3 2
13 3 0 2 3 0 2 0 3 0 2 3 0 0
14 3 0 3 0 2 1 0 1 3 3 3 0 1 3
9 3 1 1 3 0 3 0 2 3
5 3 3 1 3 3
5 3 0 2 3 0
14 3 0 3 1 3 1 2 0 1 1 3 0 0 0
2 3 3
2 3 3
9 3 1 1 1 1 1 1 0 1
10 3 3 1 3 3 3 0 0 1 3
5 3 1 3 3 2
6 3 1 3 0 0 0
1 3
1 3
7 3 1 0 3 3 3 3
4 3 0 3 3
8 3 0 3 1 3 0 2 3
4 3 0 3 3
13 3 0 0 2 1 3 0 1 1 1 1 1 1
6 3 0 2 3 1 1
1 3
8 3 0 3 1 2 0 3 0
19 3 3 0 1 1 1 2 1 3 1 3 3 0 2 0 1 3 1 0
8 3 0 3 3 0 1 2 3
3 3 0 3
2 3 3
9 3 3 0 0 0 3 0 0 1
9 3 3 0 2 3 2 3 0 3
4 3 2 0 3
12 3 0 1 3 3 0 1 3 3 0 3 0
3 3 3 0
12 3 0 1 3 3 0 1 0 3 3 1 3
6 3 2 0 1 1 3
6 3 0 3 1 2 0
2 3 3
13 3 0 3 1 3 3 1 3 3 3 0 1 0
3 3 1 2
27 3 0 2 3 1 1 1 2 0 3 0 3 0 2 1 1 2 3 1 1 3 1 1 1 2 0 3
4 3 0 3 3
3 3 3 0
4 3 1 2 3
6 3 1 3 1 3 3
7 3 3 2 3 0 1 1
1 3
7 3 3 2 3 0 3 0
10 3 3 3 0 2 0 3 1 2 3
4 3 3 1 3
11 3 3 1 1 1 1 1 3 3 1 1
1 3
7 3 3 3 1 1 3 0
16 3 0 0 2 1 1 2 0 3 3 0 2 1 3 3 2
11 3 0 3 0 2 3 3 0 0 3 0
1 3
1 3
7 3 0 3 3 1 0 0
2 3 3
2 3 3
16 3 0 3 0 1 3 3 0 1 0 2 1 1 1 3 0
2 3 3
7 3 0 3 1 3 1 3
7 3 1 0 3 3 1 0
20 3 3 1 3 3 0 3 0 0 2 3 1 1 3 3 3 3 3 3 0
12 3 0 3 0 1 3 3 0 2 3 0 3
12 3 1 3 0 2 2 0 3 0 2 0 3
17 3 0 3 1 2 2 0 3 1 2 1 1 1 2 0 2 3
1 3
11 3 1 3 1 3 3 0 1 3 3 0
3 3 1 2
2 3 3
1 3
6 3 3 1 1 0 3
6 3 2 0 3 0 0
8 3 3 0 1 1 1 1 3
3 3 3 0
5 3 3 1 0 2
2 3 3
2 3 0
9 3 0 2 3 0 2 0 3 2
14 3 3 1 1 1 1 1 1 3 3 2 0 3 0
3 3 3 0
1 3
12 3 3 0 2 2 0 3 0 2 0 3 0
10 3 0 3 0 2 2 2 3 0 0
2 3 3
16 3 1 1 1 1 3 0 3 3 0 3 0 1 2 0 3
13 3 3 0 2 1 1 1 1 2 0 2 3 2
3 3 1 3
10 3 0 2 3 1 3 3 0 3 3
4 3 0 3 0
16 3 0 3 0 2 3 0 0 3 3 1 3 0 3 1 3
11 3 1 0 3 3 3 0 1 1 1 0
10 3 3 2 0 2 1 1 1 1 2
2 3 3
14 3 0 3 3 1 3 3 0 1 2 0 3 0 1
5 3 0 2 1 3
3 3 1 3
6 3 0 3 1 3 0
3 3 3 2
2 3 0
13 3 1 3 2 0 2 0 1 2 1 1 3 1
10 3 0 3 1 1 1 1 3 1 3
7 3 3 1 2 0 3 0
4 3 0 2 3
7 3 0 3 1 2 1 0
4 3 0 3 3
16 3 0 3 0 0 3 0 3 1 3 3 1 2 0 1 3
4 3 0 3 0
3 3 3 0
9 3 0 3 1 2 1 2 1 3
8 3 2 0 3 0 0 1 3
1 3
36 3 0 3 0 2 0 0 1 1 3 3 1 3 3 0 0 3 0 0 3 0 1 3 3 0 3 3 0 0 1 3 0 1 2 3 0
11 3 1 3 0 2 0 3 0 3 0 3
10 3 0 3 1 3 3 0 1 3 2
3 3 3 0
12 3 3 0 2 3 1 3 3 3 1 3 0
20 3 3 0 1 1 1 1 1 0 2 0 3 1 2 3 0 2 1 3 0
4 3 1 3 0
17 3 3 0 2 0 3 0 1 3 3 0 1 3 3 3 0 2
6 3 0 1 0 1 3
3 3 3 2
2 3 3
5 3 0 3 0 0
6 3 0 3 1 3 3
11 3 1 3 0 1 1 2 3 2 3 2
10 3 3 1 3 3 1 2 1 1 3
5 3 3 1 3 3
8 3 0 2 3 0 0 1 3
7 3 0 3 3 1 0 0
7 3 2 1 2 1 3 2
3 3 0 3
1 3
5 3 0 2 3 0
6 3 0 3 0 1 2
4 3 0 3 3
7 3 3 1 3 3 3 3
12 3 0 3 0 3 1 3 0 1 2 3 2
1 3
7 3 0 2 3 0 0 3
12 3 1 3 0 0 3 3 1 0 1 3 3
19 3 3 3 0 2 1 3 0 0 0 3 3 3 1 3 0 3 3 0
3 3 0 3
17 3 0 3 0 1 2 3 0 3 1 3 3 0 1 1 2 3
13 3 3 1 3 3 0 3 0 2 0 1 3 0
11 3 0 2 3 0 2 0 3 1 2 3
4 3 0 3 3
3 3 3 0
1 3
8 3 0 3 1 3 2 0 3
9 3 3 0 0 3 3 2 0 2
8 3 3 0 2 1 3 1 3
10 3 0 2 3 0 2 1 1 3 3
11 3 0 3 0 1 3 3 3 2 0 0
10 3 3 0 1 0 0 3 3 1 1
6 3 0 3 0 2 3
8 3 0 1 3 3 0 2 0
10 3 3 0 2 0 3 1 0 2 3
4 3 0 3 0
2 3 0
9 3 0 3 1 3 3 0 0 0
4 3 0 2 0
13 3 3 2 3 0 3 1 2 0 3 0 0 0
13 3 3 0 1 1 3 2 0 1 1 3 0 0
4 3 0 2 3
4 3 0 3 0
3 3 0 3
4 3 3 0 0
3 3 0 3
5 3 0 3 0 3
19 3 3 0 1 1 1 1 2 0 3 2 0 3 0 1 1 1 0 1
23 3 0 3 1 2 0 1 3 1 3 3 0 1 2 0 3 0 2 0 3 0 3 3
3 3 3 0
2 3 3
20 3 3 0 3 3 1 0 2 2 0 3 0 1 3 3 2 1 2 0 3
4 3 1 3 0
15 3 1 3 0 2 0 3 1 2 1 2 0 3 3 0
3 3 0 3
7 3 1 3 0 1 1 3
2 3 3
25 3 2 2 3 1 2 0 1 3 3 1 2 1 1 1 2 0 3 2 2 1 1 2 2 0
3 3 0 3
7 3 3 3 0 2 0 3
17 3 3 2 0 3 0 2 3 1 3 3 1 3 1 1 3 0
3 3 0 2
2 3 3
3 3 0 3
3 3 2 2
7 3 0 3 0 3 0 3
13 3 3 2 3 3 1 3 3 3 1 3 0 2
8 3 0 3 3 2 3 0 1
5 3 0 3 1 0
2 3 3
2 3 3
2 3 2
2 3 3
17 3 0 1 1 1 1 2 0 3 1 2 0 1 2 0 1 3
6 3 3 0 1 0 1
7 3 0 3 3 1 3 3
2 3 3
4 3 0 2 3
13 3 0 2 1 3 1 3 3 0 2 1 3 0
9 3 0 3 1 2 0 3 3 3
12 3 1 3 0 2 0 3 0 2 3 0 1
14 3 0 3 0 1 1 1 1 0 0 1 3 3 3
2 3 3
2 3 3
6 3 3 1 3 3 3
25 3 1 2 0 1 1 1 2 1 3 0 2 0 1 3 3 0 3 3 0 2 0 1 3 3
3 3 0 3
14 3 0 3 1 2 0 3 0 1 1 2 3 1 0
8 3 0 3 1 2 3 0 2
16 3 3 1 3 3 0 0 2 3 0 1 1 3 2 1 0
7 3 0 3 0 1 2 3
9 3 0 0 0 3 1 3 3 0
3 3 0 3
3 3 1 3
16 3 0 2 1 3 0 1 1 3 0 1 1 3 1 2 3
4 3 3 0 2
12 3 0 3 1 0 2 0 0 2 0 3 0
3 3 0 3
6 3 0 3 2 0 3
6 3 0 3 0 2 0
3 3 1 3
4 3 3 2 0
2 3 3
25 3 3 1 3 3 1 1 1 1 1 3 0 1 2 3 3 2 3 0 2 0 3 0 1 2
4 3 0 2 3
3 3 1 3
4 3 0 3 0
3 3 1 3
7 3 0 2 3 0 2 3
7 3 1 3 1 3 3 3
2 3 3
1 3
3 3 1 3
10 3 3 1 3 3 0 0 3 2 3
33 3 1 3 1 1 1 0 3 0 1 3 3 0 1 3 3 0 1 3 3 0 1 3 3 1 2 2 0 3 0 2 0 0
1 3
2 3 0
5 3 0 3 3 0
4 3 0 3 3
3 3 0 3
1 3
4 3 0 2 3
30 3 0 3 0 3 1 2 0 3 1 0 2 2 2 3 1 3 3 1 3 0 1 3 0 2 3 0 0 1 3
3 3 3 0
8 3 0 3 0 1 3 3 3
10 3 0 3 0 2 0 0 0 3 0
13 3 0 3 0 3 1 2 2 3 1 3 3 2
2 3 3
8 3 0 2 3 0 2 1 2
9 3 0 3 1 2 2 3 1 3
3 3 1 3
13 3 3 0 2 3 3 0 2 0 3 0 1 2
8 3 3 0 2 1 0 0 1
8 3 3 1 0 0 0 0 3
9 3 0 3 0 2 0 3 0 2
12 3 3 1 3 3 3 0 3 0 1 2 3
16 3 0 1 2 0 3 0 1 3 3 0 3 2 0 1 3
1 3
7 3 3 0 0 1 3 0
1 3
3 3 1 3
15 3 0 3 1 3 3 1 3 3 1 3 0 2 0 1
11 3 1 3 0 2 0 1 3 3 3 0
2 3 3
5 3 1 3 2 3
7 3 0 3 1 3 0 2
2 3 3
4 3 0 2 3
8 3 3 0 2 0 3 0 1
5 3 1 3 2 3
4 3 3 0 1
2 3 3
7 3 3 1 1 3 2 0
7 3 0 3 0 3 1 3
8 3 0 3 1 2 2 0 1
2 3 3
3 3 3 3
5 3 3 0 0 0
8 3 3 1 2 1 1 1 0
4 3 0 2 3
3 3 1 3
10 3 0 1 3 3 1 2 2 0 3
4 3 3 3 2
18 3 0 3 0 1 3 3 3 0 2 1 2 0 2 1 2 1 3
12 3 2 0 0 3 0 1 0 2 0 2 0
8 3 0 3 3 1 3 2 2
3 3 0 3
2 3 1
18 3 1 3 1 3 3 0 1 3 3 0 3 1 3 3 0 2 1
3 3 1 3
12 3 3 0 1 2 1 3 1 3 2 0 3
6 3 0 3 3 0 0
3 3 3 2
5 3 1 1 3 0
6 3 2 0 3 0 2
6 3 0 2 3 0 2
2 3 3
3 3 3 2
2 3 3
2 3 2
2 3 3
5 3 3 0 0 3
6 3 0 1 2 1 3
6 3 3 1 3 3 3
2 3 3
4 3 0 3 0
13 3 3 1 1 2 0 2 3 3 3 3 3 0
6 3 3 0 2 0 2
3 3 0 3
9 3 3 2 0 2 0 3 0 2
2 3 3
11 3 0 3 1 0 1 3 3 1 3 0
12 3 3 2 0 2 0 3 0 1 3 3 0
3 3 0 3
3 3 3 0
10 3 0 2 0 1 0 1 3 3 1
3 3 1 3
12 3 0 3 3 0 0 1 3 0 1 1 3
11 3 1 3 1 3 3 3 1 1 1 3
19 3 0 3 0 1 1 3 3 0 3 1 0 1 3 3 1 1 3 0
11 3 1 3 0 2 1 3 1 3 3 3
14 3 1 3 0 2 0 3 0 1 2 3 0 3 0
3 3 3 0
1 3
13 3 3 1 3 3 1 2 1 1 2 1 3 1
1 3
7 3 3 0 3 3 1 2
27 3 0 3 0 1 2 1 3 2 1 1 1 2 0 3 0 3 1 0 1 3 3 1 3 0 0 0
8 3 0 3 1 2 1 0 1
3 3 0 2
17 3 3 1 3 3 3 1 0 0 2 0 3 0 2 2 2 3
2 3 3
3 3 3 0
18 3 1 1 3 3 0 1 0 1 3 0 2 0 3 1 2 1 0
3 3 3 2
14 3 1 3 0 2 2 2 1 0 1 0 2 1 0
3 3 3 0
4 3 3 1 2
13 3 0 3 1 3 1 3 0 1 2 1 3 0
14 3 1 3 2 0 1 2 3 0 2 3 1 3 3
7 3 3 2 0 0 1 1
10 3 1 3 1 3 2 2 0 3 0
5 3 0 3 0 1
4 3 0 2 3
1 3
4 3 0 2 3
13 3 0 3 0 1 3 3 3 2 0 0 1 3
2 3 0
17 3 3 1 3 3 0 3 1 2 1 1 0 2 1 1 3 3
8 3 0 3 1 3 0 2 3
3 3 2 2
6 3 1 1 0 3 1
5 3 3 0 1 3
10 3 3 1 3 3 3 1 3 3 3
6 3 3 0 0 1 3
2 3 3
3 3 1 3
7 3 0 2 3 0 1 3
2 3 1
6 3 3 1 3 3 3
2 3 3
6 3 0 3 0 1 0
14 3 0 3 0 3 3 1 1 3 2 1 2 0 3
2 3 1
8 3 1 1 3 1 3 3 3
3 3 0 3
3 3 3 0
5 3 0 3 0 2
2 3 3
13 3 3 0 0 3 3 3 3 3 0 1 0 3
6 3 0 3 1 3 3
5 3 3 0 0 0
17 3 0 3 1 3 0 3 0 1 2 1 3 3 3 0 1 3
6 3 3 3 0 0 0
3 3 0 3
8 3 3 1 3 3 1 3 3
5 3 2 0 1 3
7 3 3 0 1 1 3 1
12 3 0 3 0 1 1 1 1 1 3 0 3
11 3 0 3 0 2 0 1 2 0 3 0
3 3 1 3
13 3 3 0 0 3 0 0 0 3 3 1 2 1
15 3 3 1 3 3 3 1 0 3 1 3 3 3 0 3
3 3 3 0
8 3 0 3 3 2 3 1 0
3 3 1 3
8 3 0 1 2 2 3 1 0
3 3 0 3
4 3 0 2 3
2 3 3
6 3 3 0 0 0 1
2 3 3
3 3 2 2
1 3
25 3 3 0 1 0 1 3 3 3 0 3 1 3 0 2 0 1 0 1 1 3 0 1 0 0
15 3 0 3 1 3 0 3 0 1 1 3 3 0 2 0
3 3 1 3
23 3 3 0 0 1 2 2 0 3 0 2 1 3 0 2 0 3 1 2 0 3 1 0
7 3 3 1 1 3 2 0
1 3
2 3 0
2 3 3
1 3
18 3 0 3 0 1 2 0 3 0 3 0 0 3 1 3 0 2 3
3 3 3 0
11 3 3 1 1 1 1 0 0 3 1 3
2 3 3
2 3 3
2 3 3
10 3 0 3 3 0 2 1 1 3 3
2 3 0
3 3 1 3
15 3 0 3 0 3 1 3 0 3 0 1 3 3 0 3
2 3 3
6 3 0 1 2 0 3
6 3 3 0 2 1 3
2 3 3
3 3 0 2
16 3 3 2 0 2 3 1 3 0 2 1 0 0 2 3 0
10 3 1 3 1 1 1 3 3 2 2
5 3 3 0 0 0
4 3 0 3 0
36 3 3 1 3 1 3 0 0 0 2 0 3 1 2 3 0 1 1 2 0 3 1 1 3 3 0 2 3 1 2 3 1 2 3 3 0
7 3 0 3 0 1 3 3
8 3 3 1 0 1 3 3 3
6 3 1 3 1 3 3
2 3 3
4 3 3 0 2
18 3 3 2 0 2 0 1 3 1 0 1 3 0 0 1 3 0 0
1 3
9 3 3 0 1 1 1 1 2 0
2 3 3
16 3 3 0 2 0 3 0 1 1 3 1 3 0 2 3 1
4 3 3 0 2
5 3 0 2 3 0
5 3 0 3 3 0
5 3 0 1 2 1
6 3 1 1 3 3 1
10 3 3 0 1 1 1 1 1 2 3
5 3 3 2 0 0
5 3 0 2 3 0
6 3 0 3 0 1 2
3 3 3 0
2 3 3
11 3 1 1 1 1 1 3 3 2 1 0
15 3 3 0 2 1 0 3 3 2 0 3 0 1 2 3
11 3 0 3 0 3 0 3 3 0 1 0
10 3 0 3 0 1 3 3 3 0 2
6 3 0 3 0 2 1
3 3 3 2
10 3 2 0 3 0 2 2 0 3 0
3 3 3 2
1 3
9 3 0 3 0 3 1 0 3 2
5 3 3 3 0 1
2 3 3
1 3
2 3 3
14 3 3 0 2 1 3 0 1 2 0 2 3 1 2
4 3 0 3 0
2 3 3
11 3 3 0 1 2 3 0 1 3 3 3
7 3 3 1 3 3 3 0
3 3 0 0
21 3 0 3 1 2 1 1 1 1 1 2 1 3 0 2 1 1 3 1 1 3
16 3 0 1 3 3 3 3 3 3 2 0 0 0 1 2 2
2 3 3
4 3 0 3 0
8 3 1 3 1 3 3 0 2
4 3 3 3 0
5 3 1 1 2 3
3 3 1 3
6 3 1 0 3 3 3
4 3 0 2 3
2 3 3
3 3 0 1
7 3 1 3 0 0 1 3
1 3
8 3 0 3 3 0 0 1 3
7 3 0 3 0 3 3 0
21 3 0 3 0 1 3 1 3 3 1 0 1 3 3 3 1 3 1 3 3 3
6 3 0 3 0 3 3
2 3 0
4 3 0 2 3
6 3 1 3 0 0 0
31 3 3 0 2 1 1 3 1 1 2 3 0 1 3 3 3 0 1 1 2 0 2 3 0 2 0 3 0 1 3 3
3 3 1 3
9 3 0 3 0 3 1 3 0 3
2 3 3
6 3 0 3 0 2 3
4 3 0 1 2
2 3 3
2 3 3
1 3
4 3 0 3 0
10 3 3 1 3 3 3 0 2 3 0
2 3 1
8 3 0 1 3 3 1 2 3
4 3 1 3 0
2 3 3
14 3 0 3 0 2 2 0 0 3 3 3 3 3 3
12 3 3 0 2 1 3 1 3 3 3 2 3
12 3 3 0 1 1 1 2 0 3 1 0 2
10 3 3 0 0 2 3 1 2 3 0
5 3 3 1 3 3
4 3 3 1 2
13 3 0 3 1 2 2 0 3 1 3 0 1 2
4 3 0 2 3
10 3 0 2 3 0 0 1 3 0 2
10 3 1 3 1 3 0 3 0 3 0
8 3 0 3 0 3 3 0 0
4 3 3 0 0
9 3 3 1 1 3 1 3 0 2
17 3 3 0 1 1 0 3 1 0 1 3 0 1 1 1 0 2
4 3 3 1 3
12 3 0 3 1 2 0 3 1 1 2 0 3
5 3 0 3 3 0
6 3 3 0 2 1 2
2 3 3
17 3 3 0 1 3 2 0 1 3 1 1 0 2 1 1 0 2
8 3 2 0 3 0 0 0 1
13 3 1 1 3 1 3 3 3 0 2 2 0 3
4 3 3 1 3
2 3 3
2 3 3
4 3 3 0 2
7 3 3 1 2 1 3 0
7 3 0 3 0 2 1 3
4 3 0 2 3
9 3 0 3 0 1 2 0 3 0
13 3 1 3 1 3 0 2 1 2 0 3 1 2
21 3 0 3 1 3 0 2 3 0 3 1 3 3 0 1 3 3 0 3 0 3
4 3 3 0 0
4 3 0 3 3
1 3
19 3 0 3 3 0 1 3 1 1 0 1 3 3 1 2 1 1 1 1
1 3
3 3 0 3
3 3 0 3
3 3 0 3
4 3 2 0 3
15 3 0 3 0 0 1 2 2 3 1 3 3 3 0 0
2 3 1
9 3 0 3 0 3 1 2 1 3
28 3 3 3 1 3 3 0 1 2 0 3 0 1 3 3 0 3 0 3 1 2 1 1 1 3 2 1 3
3 3 0 3
2 3 3
4 3 0 3 3
3 3 1 3
9 3 0 3 1 0 1 3 3 0
16 3 1 3 0 1 1 3 2 3 0 1 3 1 0 3 3
2 3 3
5 3 1 3 2 3
7 3 3 1 2 3 0 3
3 3 3 0
3 3 1 3
7 3 0 3 1 2 0 3
9 3 3 1 3 3 1 3 3 0
1 3
4 3 3 0 3
1 3
13 3 3 1 2 1 1 2 0 3 3 0 0 0
14 3 1 3 1 1 1 3 1 3 0 0 0 3 0
12 3 3 0 2 1 1 3 0 0 3 3 0
4 3 0 3 2
3 3 0 3
3 3 3 0
8 3 3 2 2 2 3 0 0
7 3 0 3 1 0 1 0
6 3 0 3 1 0 0
3 3 3 0
9 3 0 3 0 0 1 2 3 0
2 3 3
8 3 0 2 2 1 1 1 0
6 3 3 1 2 3 0
5 3 3 1 1 1
20 3 1 3 0 3 3 2 3 0 0 2 3 1 1 1 1 1 1 3 0
6 3 1 1 3 0 2
20 3 0 3 0 1 3 3 0 2 0 3 3 1 2 2 3 1 0 2 3
12 3 0 3 0 3 2 3 1 1 2 3 3
9 3 0 3 3 0 0 1 1 3
2 3 3
3 3 3 2
7 3 0 3 1 2 3 0
12 3 0 3 1 0 1 3 3 0 3 1 3
4 3 0 1 2
2 3 0
7 3 1 3 0 2 1 2
7 3 0 2 3 0 1 3
3 3 1 3
3 3 0 0
1 3
5 3 0 1 0 0
5 3 3 1 3 3
3 3 0 3
7 3 0 3 0 2 3 0
3 3 3 3
10 3 0 1 0 3 0 0 2 0 3
8 3 0 3 1 2 1 2 3
24 3 3 2 0 0 0 0 3 3 3 1 1 3 1 1 1 3 1 3 0 2 3 1 2
3 3 3 0
4 3 3 1 0
2 3 3
3 3 3 0
21 3 3 0 1 1 2 3 1 0 1 3 3 0 3 0 1 2 2 0 2 3
5 3 2 0 3 0
4 3 3 2 1
32 3 3 1 3 3 1 1 3 1 1 3 1 3 1 0 0 3 3 3 1 0 2 0 1 2 1 1 2 0 3 0 0
22 3 3 0 1 0 1 3 3 3 3 1 0 2 0 3 1 0 1 3 3 0 3
16 3 0 2 0 0 2 0 3 0 1 2 3 1 3 3 3
7 3 3 1 2 0 0 3
7 3 2 0 3 0 0 0
10 3 3 0 1 3 1 3 3 3 3
8 3 3 3 1 3 3 3 2
15 3 1 3 0 0 3 3 0 1 1 3 3 0 3 3
8 3 0 3 1 2 0 1 3
10 3 1 0 3 0 0 1 3 3 3
12 3 0 2 1 3 1 3 3 1 2 1 3
6 3 0 3 0 1 0
5 3 3 2 0 0
39 3 0 3 3 1 3 3 1 3 3 0 1 3 2 2 3 1 3 3 1 2 1 3 0 1 1 2 3 0 1 0 2 3 1 2 0 2 1 3
3 3 3 0
10 3 0 3 0 3 0 2 2 1 1
1 3
16 3 3 1 3 3 0 3 0 3 0 1 0 2 3 0 2
2 3 0
4 3 0 3 3
10 3 0 3 1 3 0 1 2 1 3
32 3 0 3 0 1 3 3 0 3 3 3 0 0 3 3 0 1 1 3 3 1 3 0 0 1 3 0 1 1 1 1 0
6 3 1 2 0 1 3
13 3 3 1 3 3 1 0 3 3 2 0 0 3
27 3 0 3 0 0 2 1 0 1 1 3 3 0 1 0 2 3 0 3 1 2 3 0 1 1 1 3
3 3 0 3
5 3 0 3 1 3
3 3 1 3
8 3 0 3 0 3 1 2 1
3 3 0 3
12 3 0 3 1 3 1 3 3 0 3 1 3
27 3 1 3 2 0 0 3 3 0 0 3 0 1 0 1 3 3 1 3 0 2 0 3 0 1 0 0
17 3 3 0 1 1 1 1 1 2 0 3 0 2 3 2 0 3
13 3 3 0 0 3 3 1 3 3 0 2 0 3
5 3 1 0 1 3
11 3 0 3 0 3 0 2 0 3 0 2
4 3 1 1 3
12 3 3 0 2 3 1 3 1 3 2 0 3
14 3 0 3 0 1 3 1 2 2 0 3 0 0 3
4 3 0 3 3
5 3 3 1 3 3
25 3 0 3 1 3 0 3 0 3 0 1 1 3 2 0 3 1 3 3 1 2 1 3 1 1
13 3 0 3 1 2 2 3 2 0 0 1 1 3
5 3 1 1 3 0
4 3 3 0 0
4 3 0 1 0
9 3 3 1 3 3 3 3 3 0
4 3 3 0 0
12 3 0 3 1 0 1 3 3 3 1 3 0
2 3 3
9 3 0 3 0 1 3 3 1 3
7 3 0 3 1 3 1 2
1 3
3 3 3 2
3 3 0 3
15 3 3 0 1 1 1 0 1 3 3 3 0 3 1 3
3 3 0 1
10 3 2 0 3 0 1 1 1 2 3
1 3
12 3 1 3 0 1 3 3 3 3 0 2 1
8 3 0 3 0 1 3 3 3
1 3
4 3 0 2 3
2 3 0
12 3 1 1 1 3 1 1 1 1 1 1 3
15 3 3 1 3 0 3 3 3 3 0 0 1 0 3 1
3 3 1 3
2 3 1
6 3 1 1 3 3 3
2 3 3
10 3 3 3 0 1 1 1 2 3 2
3 3 3 0
10 3 1 3 3 2 0 1 1 1 1
3 3 3 2
12 3 0 1 3 3 1 0 1 2 0 0 3
5 3 3 1 2 3
3 3 0 3
10 3 0 1 2 1 2 3 0 0 3
13 3 3 0 3 3 0 3 0 1 1 3 0 3
12 3 0 3 0 0 3 0 1 3 3 0 2
4 3 3 3 2
5 3 1 1 1 2
4 3 3 2 3
2 3 3
5 3 0 3 3 0
3 3 2 1
15 3 1 3 1 3 3 0 1 3 3 0 3 1 3 1
4 3 0 1 2
2 3 3
3 3 1 2
20 3 1 3 0 1 3 3 3 3 0 0 3 0 1 1 1 2 1 0 0
9 3 0 3 0 3 1 3 1 3
6 3 0 3 1 3 3
2 3 3
3 3 1 3
3 3 3 2
12 3 0 2 3 0 1 2 0 1 0 3 0
4 3 3 3 2
6 3 0 3 3 0 0
2 3 0
7 3 0 3 1 2 0 3
4 3 1 1 3
9 3 0 3 3 3 0 2 0 3
3 3 1 3
8 3 0 3 0 3 3 0 2
2 3 3
2 3 3
2 3 3
17 3 0 1 1 3 3 3 1 0 2 0 1 2 1 2 0 3
4 3 0 3 0
3 3 3 0
4 3 0 2 3
6 3 3 1 0 3 1
3 3 0 3
15 3 3 1 3 3 1 1 3 2 0 3 0 0 1 3
5 3 0 3 0 2
4 3 1 0 0
2 3 3
10 3 3 0 2 0 3 1 2 1 3
3 3 1 1
12 3 1 3 0 0 1 1 3 0 2 0 3
16 3 3 1 1 1 3 0 0 1 1 1 2 3 1 3 3
8 3 0 3 3 0 0 1 3
11 3 2 0 3 0 1 2 0 3 0 1
9 3 0 1 3 3 0 1 1 3
3 3 3 0
1 3
10 3 0 3 1 2 1 1 2 0 3
5 3 0 2 3 0
3 3 1 3
5 3 0 3 3 0
9 3 0 3 0 1 3 3 3 2
17 3 3 1 3 3 0 0 3 1 2 3 1 2 1 1 3 0
3 3 3 0
4 3 3 0 1
4 3 0 1 0
2 3 0
1 3
9 3 0 3 1 2 2 0 3 3
8 3 3 0 0 3 3 3 0
6 3 3 0 2 0 3
15 3 0 3 1 3 3 2 1 3 3 0 1 2 0 3
3 3 3 0
10 3 2 0 3 0 2 3 1 3 1
15 3 0 0 2 3 0 2 0 3 1 0 2 3 0 3
3 3 1 3
3 3 0 3
19 3 0 2 0 3 1 3 3 3 1 3 3 1 2 2 3 2 0 0
5 3 3 0 0 0
12 3 0 3 0 2 0 0 1 2 0 2 3
2 3 3
3 3 3 1
5 3 0 2 0 0
1 3
8 3 3 2 2 2 1 3 1
9 3 3 0 0 0 3 3 3 3
2 3 3
6 3 0 2 1 3 0
2 3 3
3 3 1 3
1 3
2 3 3
10 3 0 3 3 1 3 3 1 3 3
3 3 1 3
8 3 0 3 0 1 3 3 3
1 3
6 3 0 1 2 0 2
8 3 0 3 3 2 1 1 3
18 3 3 0 2 1 1 3 3 1 2 2 0 3 0 1 0 3 1
3 3 0 1
4 3 0 3 3
28 3 0 3 1 2 0 0 0 3 3 3 0 1 2 1 1 1 2 3 2 0 2 1 1 1 3 3 3
4 3 0 3 3
9 3 0 3 0 1 3 3 3 0
1 3
14 3 0 3 1 3 3 0 2 2 0 1 1 3 0
3 3 0 3
15 3 1 0 3 3 0 3 0 0 3 0 1 0 1 2
3 3 0 1
18 3 3 3 0 3 3 0 2 1 3 0 0 1 1 1 1 3 0
3 3 2 2
3 3 0 1
5 3 1 3 0 2
8 3 0 3 1 1 3 3 1
2 3 0
1 3
3 3 0 3
4 3 0 3 0
6 3 3 1 3 3 0
19 3 3 0 1 3 2 1 2 0 3 0 2 0 3 1 3 3 3 0
14 3 0 1 2 3 1 3 3 1 0 1 2 1 0
10 3 0 3 1 2 3 0 2 1 3
1 3
8 3 0 3 0 1 0 1 3
7 3 3 2 0 0 1 3
11 3 0 3 0 0 0 1 3 3 3 2
5 3 3 3 0 3
3 3 3 0
5 3 0 3 1 0
2 3 3
2 3 3
17 3 0 3 1 0 1 2 1 2 0 3 0 1 1 3 0 3
15 3 0 1 3 3 0 3 0 0 1 3 3 3 2 0
2 3 3
6 3 3 1 3 3 3
8 3 0 2 1 1 3 0 2
2 3 3
4 3 0 3 0
8 3 1 1 3 1 3 3 3
6 3 3 1 3 3 3
5 3 3 1 2 1
2 3 3
5 3 1 1 1 3
10 3 3 0 1 1 2 0 3 3 3
3 3 3 0
6 3 0 1 2 1 3
1 3
7 3 0 3 0 1 2 0
11 3 0 3 1 3 0 1 2 0 3 0
5 3 0 2 3 2
8 3 0 3 0 2 3 1 3
6 3 0 3 0 2 3
6 3 0 0 3 3 3
3 3 3 2
10 3 3 2 1 1 3 0 3 3 2
25 3 0 2 3 1 0 0 1 3 3 3 1 3 0 2 0 3 1 3 0 3 1 3 3 0
5 3 3 3 3 0
2 3 3
2 3 0
14 3 3 1 3 3 0 3 1 3 1 3 0 0 0
3 3 0 3
9 3 0 3 0 3 0 1 2 3
6 3 1 3 0 0 3
6 3 1 1 1 3 0
18 3 0 3 1 0 1 3 3 0 2 3 1 3 3 0 1 0 0
2 3 3
5 3 3 0 0 3
13 3 3 2 1 3 0 3 0 3 0 3 3 0
4 3 3 0 0
24 3 1 3 0 2 1 2 1 1 3 0 3 1 2 1 3 0 1 3 3 3 1 3 3
6 3 0 3 3 1 2
6 3 2 0 1 1 3
1 3
5 3 0 1 3 3
3 3 0 3
3 3 0 3
21 3 1 3 0 2 0 3 0 3 1 0 1 2 1 3 0 2 2 0 3 0
16 3 1 3 1 3 3 3 0 3 1 1 2 0 3 3 3
7 3 0 1 1 1 1 1
22 3 0 3 1 3 2 0 1 3 0 0 1 3 0 2 0 3 3 0 1 1 3
4 3 1 1 2
8 3 0 3 1 2 1 3 0
27 3 2 0 3 0 2 0 3 0 3 0 1 3 3 0 2 1 3 2 0 2 0 3 1 2 0 0
3 3 0 3
3 3 0 3
3 3 3 0
9 3 0 3 1 0 0 1 2 3
3 3 0 3
2 3 3
3 3 1 3
15 3 0 2 3 3 0 1 3 3 3 2 0 1 3 0
1 3
6 3 3 1 3 3 3
3 3 0 3
1 3
8 3 0 3 1 3 1 1 1
2 3 3
9 3 3 1 2 3 0 2 3 0
3 3 0 3
4 3 1 3 0
5 3 1 3 1 3
12 3 0 3 1 1 3 0 0 1 2 0 3
1 3
1 3
14 3 1 2 2 1 2 1 1 1 3 0 0 1 3
2 3 3
3 3 1 3
5 3 1 3 0 1
19 3 0 3 0 2 0 1 2 2 0 3 3 0 1 2 0 3 1 3
2 3 3
2 3 3
2 3 3
16 3 3 0 2 0 3 1 3 0 1 1 1 1 1 1 0
3 3 0 3
7 3 2 3 0 2 0 0
2 3 3
5 3 1 0 0 0
3 3 2 3
1 3
11 3 0 3 3 2 1 0 1 3 3 3
3 3 0 3
4 3 3 0 2
6 3 0 3 0 3 0
8 3 3 1 3 3 3 2 1
8 3 0 3 0 1 2 1 3
1 3
6 3 0 2 3 0 2
1 3
14 3 1 1 1 3 1 2 0 2 0 1 3 3 3
2 3 0
11 3 0 3 3 1 3 3 1 2 1 0
14 3 3 1 0 0 3 0 1 2 2 0 3 0 2
5 3 2 0 3 0
9 3 0 3 1 2 2 0 2 3
10 3 0 3 1 2 1 1 2 0 3
31 3 1 3 0 1 1 1 3 3 0 3 3 3 3 0 1 3 3 0 3 1 2 1 2 0 2 3 0 0 1 3
7 3 0 3 1 2 0 3
4 3 1 3 0
5 3 3 3 3 3
4 3 0 3 3
1 3
5 3 3 1 3 3
2 3 0
4 3 0 3 0
3 3 1 3
10 3 3 1 3 3 0 2 1 1 2
2 3 0
7 3 0 3 0 1 0 0
2 3 3
14 3 3 1 2 1 1 2 3 2 0 2 1 3 0
4 3 0 2 3
5 3 0 1 0 0
3 3 0 2
13 3 0 3 0 1 0 1 2 1 3 0 1 3
5 3 3 0 1 0
19 3 0 3 1 3 1 1 1 1 1 1 3 1 3 0 1 1 1 2
7 3 0 3 3 1 3 3
4 3 3 3 2
10 3 3 0 2 1 3 0 3 3 0
25 3 0 1 1 3 2 1 1 0 1 3 3 3 3 0 0 0 1 1 3 1 3 3 0 0
2 3 3
7 3 3 1 3 0 3 3
3 3 0 3
5 3 0 3 0 0
2 3 3
7 3 1 3 0 1 2 3
3 3 0 3
16 3 2 0 3 0 1 1 1 1 1 1 1 1 1 1 3
5 3 0 2 3 0
1 3
10 3 3 1 3 0 3 0 3 3 2
3 3 1 3
15 3 0 2 1 1 3 0 0 1 3 0 2 0 3 0
11 3 3 1 3 3 1 1 3 1 1 3
2 3 3
6 3 0 3 0 2 3
1 3
11 3 0 3 1 3 3 3 1 0 1 0
13 3 1 3 1 3 1 1 1 1 1 1 0 1
9 3 0 3 1 2 1 1 0 2
4 3 0 3 3
8 3 3 0 1 1 1 1 0
1 3
22 3 1 3 3 1 3 3 1 2 2 3 3 2 3 3 1 1 3 1 3 3 0
3 3 1 3
9 3 3 0 1 1 2 3 0 2
3 3 0 3
3 3 0 3
17 3 0 3 0 1 3 3 1 0 2 2 2 3 0 2 1 2
23 3 0 3 0 1 3 3 3 0 1 0 3 1 0 1 3 3 1 1 3 3 3 0
9 3 0 3 0 1 3 3 0 3
4 3 0 3 3
3 3 1 3
5 3 3 2 0 0
25 3 3 0 1 1 1 1 1 1 3 0 1 3 3 1 1 1 1 1 1 3 0 2 0 3
2 3 3
6 3 2 2 0 1 3
4 3 0 2 3
3 3 3 0
13 3 1 3 1 3 3 1 0 2 2 1 2 3
2 3 3
1 3
3 3 0 3
5 3 1 1 3 0
11 3 0 3 0 0 1 3 3 0 3 0
9 3 3 1 3 3 0 3 1 2
4 3 0 2 3
3 3 0 3
2 3 3
4 3 3 2 1
2 3 1
2 3 0
6 3 0 3 1 2 3
13 3 0 1 0 1 1 3 1 1 1 3 1 3
4 3 1 3 0
1 3
9 3 0 3 0 3 1 3 1 3
1 3
4 3 2 0 3
2 3 3
3 3 1 3
3 3 1 3
7 3 3 0 1 1 1 0
13 3 1 3 0 2 0 3 1 3 2 0 3 0
1 3
3 3 0 3
2 3 3
3 3 0 3
12 3 1 3 0 1 2 3 1 2 2 3 2
5 3 2 0 3 0
1 3
9 3 0 3 0 3 1 3 0 2
3 3 3 3
4 3 3 0 0
6 3 0 3 0 1 0
8 3 3 0 2 0 3 1 3
8 3 3 1 3 3 3 0 2
8 3 2 3 0 1 2 3 3
7 3 0 3 0 2 3 2
3 3 0 3
1 3
5 3 0 3 0 2
2 3 0
3 3 3 0
6 3 0 3 0 2 3
2 3 3
16 3 3 1 2 3 0 1 2 0 3 1 0 1 1 3 0
1 3
6 3 3 0 1 0 2
9 3 0 3 1 0 0 1 3 3
2 3 3
13 3 0 3 1 0 1 1 3 2 1 1 0 1
4 3 0 3 3
11 3 3 0 2 3 1 3 0 1 2 3
9 3 0 3 3 1 3 3 0 3
3 3 1 3
5 3 0 3 0 3
6 3 3 1 2 1 0
2 3 3
10 3 3 1 3 3 0 3 0 3 3
11 3 0 3 0 3 1 3 3 0 1 0
7 3 0 2 3 0 2 2
1 3
10 3 3 0 2 0 3 0 2 0 3
2 3 3
4 3 0 1 0
1 3
10 3 0 3 0 0 1 1 1 1 0
5 3 0 3 0 3
4 3 1 1 3
12 3 3 0 2 0 3 1 2 2 0 2 3
8 3 3 1 0 3 3 2 1
23 3 1 0 1 3 1 2 1 2 0 3 2 0 1 3 1 3 3 0 1 1 1 2
1 3
7 3 0 1 2 3 0 3
12 3 3 1 3 3 0 2 3 0 3 0 2
6 3 3 0 1 1 3
3 3 3 0
4 3 0 2 3
7 3 0 3 1 2 3 0
1 3
5 3 3 1 2 1
13 3 3 1 3 3 0 1 2 1 0 1 3 0
5 3 1 1 3 0
2 3 3
12 3 0 1 1 3 0 3 1 2 2 0 3
8 3 0 3 1 0 1 3 3
1 3
3 3 0 3
13 3 0 3 0 3 0 1 3 3 0 3 0 0
5 3 3 2 0 0
18 3 0 3 0 0 3 0 1 2 0 1 3 1 3 3 0 3 3
4 3 1 3 2
2 3 0
18 3 3 0 1 2 0 3 3 1 3 3 3 0 0 3 3 0 1
10 3 0 3 0 1 2 0 1 1 3
12 3 0 3 1 0 1 2 3 2 0 3 0
6 3 0 3 0 1 2
1 3
11 3 0 3 1 2 3 0 1 1 1 1
1 3
22 3 3 0 2 3 0 3 3 0 0 3 0 1 2 3 0 3 1 0 1 3 3
1 3
14 3 0 2 0 1 3 3 0 3 1 2 0 3 0
2 3 1
3 3 1 3
1 3
3 3 3 0
14 3 0 3 1 0 1 3 3 0 1 3 3 1 3
2 3 3
8 3 0 3 1 2 0 3 0
42 3 0 1 3 3 1 2 2 1 3 0 0 1 1 3 1 1 1 1 1 3 1 1 1 1 1 2 0 3 1 2 0 0 1 3 3 1 2 1 3 0 0
12 3 0 3 0 3 0 0 3 1 3 1 2
4 3 0 3 0
13 3 0 3 0 3 0 0 3 3 3 1 1 3
5 3 0 2 1 3
6 3 2 0 3 0 2
7 3 0 0 3 1 3 3
20 3 3 1 3 3 1 1 3 3 1 0 1 3 3 3 0 2 0 2 3
4 3 3 0 0
11 3 0 3 0 3 0 2 0 3 2 1
32 3 0 3 1 3 1 1 1 3 0 1 0 0 1 3 3 3 0 3 0 2 0 1 3 1 1 3 0 1 3 3 0
13 3 0 3 0 1 2 3 1 3 3 0 3 3
1 3
2 3 0
3 3 3 0
3 3 0 3
13 3 0 3 3 1 3 3 0 3 0 3 0 3
8 3 0 3 1 2 0 1 3
7 3 3 0 1 1 1 3
9 3 3 0 2 0 3 0 1 0
3 3 0 3
4 3 0 2 3
9 3 0 3 0 0 3 0 2 3
6 3 0 3 0 2 3
7 3 0 3 1 3 0 3
9 3 1 3 3 1 3 3 3 0
2 3 3
11 3 0 3 1 0 2 1 1 1 1 0
4 3 3 0 2
4 3 0 3 0
8 3 2 0 3 0 2 0 2
8 3 0 3 1 0 1 0 0
10 3 0 3 1 3 3 2 0 0 0
1 3
8 3 0 3 3 3 3 0 0
16 3 1 1 3 3 3 2 0 2 1 1 3 1 3 0 0
11 3 0 3 1 3 0 3 0 3 1 3
20 3 1 3 2 0 1 3 2 3 3 1 2 1 1 1 2 0 3 0 3
13 3 1 0 0 2 0 1 2 1 1 1 1 0
4 3 3 0 2
2 3 0
3 3 0 3
6 3 0 3 1 2 3
16 3 3 3 1 3 3 1 3 3 0 1 2 1 1 3 1
11 3 0 3 1 2 3 0 2 0 0 0
6 3 0 3 0 2 0
29 3 1 3 1 3 3 0 2 0 2 0 3 0 3 1 3 3 0 1 1 1 1 3 2 3 1 3 3 0
5 3 3 0 0 0
6 3 3 2 2 2 3
4 3 1 3 0
7 3 3 0 2 1 1 1
2 3 3
9 3 0 3 0 2 1 1 0 2
9 3 0 3 1 2 0 1 1 3
2 3 3
10 3 3 0 2 0 3 0 0 1 0
3 3 0 3
7 3 3 0 2 0 3 0
3 3 1 3
3 3 0 3
2 3 3
18 3 3 3 0 1 2 0 3 1 2 1 1 1 1 1 2 0 0
3 3 3 0
7 3 0 1 2 2 0 3
2 3 3
5 3 0 0 2 3
32 3 0 1 2 1 1 3 0 1 1 1 0 1 3 1 0 2 2 2 3 0 2 1 1 1 2 0 1 2 0 3 0
12 3 3 1 3 3 0 1 3 3 3 0 2
37 3 0 3 0 1 2 0 3 0 1 1 2 0 3 0 1 3 3 0 1 3 3 3 1 0 2 0 1 3 0 3 1 2 2 3 2 3
1 3
6 3 0 3 0 2 3
22 3 1 3 0 1 2 3 0 0 3 0 1 2 1 2 1 3 0 2 0 1 2
4 3 0 2 3
2 3 2
3 3 3 0
4 3 0 2 3
4 3 1 2 1
2 3 3
13 3 3 0 0 0 2 3 3 2 0 2 3 3
2 3 3
6 3 3 0 2 0 3
14 3 3 0 0 3 3 1 3 3 3 1 2 0 2
6 3 0 3 1 2 3
9 3 0 3 3 3 1 0 3 1
2 3 0
6 3 1 1 3 0 0
3 3 0 3
9 3 3 1 3 3 3 1 3 3
3 3 3 2
1 3
7 3 3 1 3 3 3 3
7 3 0 3 0 3 0 3
2 3 3
15 3 0 3 0 1 1 3 2 0 3 0 1 2 3 2
6 3 0 2 3 0 0
13 3 0 3 0 1 1 1 1 1 1 1 3 3
8 3 1 2 1 3 1 0 0
13 3 1 1 3 3 1 2 1 2 0 3 1 3
12 3 3 2 0 0 0 0 1 2 0 3 0
2 3 0
1 3
6 3 3 0 2 0 3
9 3 0 3 3 1 3 3 3 3
12 3 0 3 0 2 0 2 3 1 3 0 1
2 3 3
2 3 3
8 3 1 3 0 1 1 1 0
34 3 3 1 3 3 1 0 2 3 1 1 3 3 3 0 1 0 1 2 1 1 2 0 3 0 1 3 3 0 0 1 3 3 3
9 3 1 1 1 1 3 1 3 0
13 3 3 1 3 3 0 3 0 1 0 3 3 3
6 3 0 2 1 3 0
11 3 1 0 3 3 1 3 1 0 3 0
11 3 0 3 0 1 2 3 0 0 0 1
8 3 0 3 0 1 3 3 0
4 3 0 3 3
5 3 0 3 1 2
24 3 1 3 0 0 1 3 0 1 2 0 3 0 1 3 3 2 0 0 3 3 1 3 3
1 3
2 3 3
2 3 3
9 3 0 3 1 0 1 2 0 3
14 3 0 3 0 2 0 3 0 1 2 0 2 3 0
4 3 1 3 0
3 3 0 3
4 3 1 1 3
8 3 0 2 3 0 0 3 3
7 3 0 3 1 2 1 0
3 3 3 0
4 3 3 0 2
3 3 0 1
20 3 0 3 0 3 3 3 3 1 3 0 3 0 1 3 3 1 3 0 0
2 3 3
5 3 3 0 0 0
6 3 0 3 1 2 3
6 3 0 3 0 1 2
3 3 0 1
7 3 0 3 0 1 3 3
5 3 0 3 1 3
14 3 3 0 1 2 0 3 1 2 1 1 3 2 2
2 3 0
4 3 3 0 0
12 3 0 3 1 2 1 1 1 2 1 3 0
3 3 0 3
3 3 0 3
6 3 1 1 3 0 1
5 3 3 0 0 0
44 3 0 1 2 1 0 3 3 1 2 1 3 3 0 3 3 3 3 0 3 0 3 1 1 1 1 3 1 3 3 0 1 3 3 2 1 3 0 2 0 3 1 0 2
23 3 0 1 3 3 0 2 3 0 2 0 3 0 2 3 3 1 3 0 2 1 1 3
1 3
5 3 0 2 1 3
2 3 3
3 3 3 3
8 3 2 0 3 0 1 1 3
1 3
3 3 0 3
3 3 0 2
5 3 0 1 2 3
16 3 0 3 0 3 3 3 0 2 0 2 0 2 0 1 0
9 3 0 3 0 2 3 1 0 3
11 3 0 1 2 0 2 3 0 1 3 3
3 3 0 2
1 3
19 3 0 3 1 0 2 2 2 3 0 0 1 3 0 0 3 3 3 0
34 3 0 3 0 1 3 3 0 1 0 3 3 0 2 3 0 3 0 1 2 0 3 0 1 3 3 0 3 3 0 1 2 3 0
1 3
14 3 3 1 1 1 2 0 3 0 0 2 0 0 2
2 3 3
11 3 0 3 1 3 3 1 3 3 3 2
6 3 0 3 1 3 3
1 3
3 3 1 3
8 3 3 0 2 0 3 0 2
2 3 3
2 3 3
8 3 0 3 3 1 3 3 3
8 3 3 3 0 2 2 1 2
7 3 3 1 3 3 1 3
7 3 0 2 2 2 0 3
3 3 0 3
4 3 0 3 0
17 3 1 1 1 0 3 0 3 0 3 2 3 2 0 1 2 3
14 3 0 1 0 1 3 3 1 3 3 0 2 3 3
8 3 3 0 0 3 3 0 3
17 3 0 0 3 0 1 1 1 1 3 3 2 2 3 1 2 3
2 3 3
2 3 1
3 3 3 3
2 3 3
4 3 0 2 3
2 3 3
1 3
6 3 0 3 1 3 0
4 3 0 0 3
10 3 0 3 0 3 1 2 1 1 0
8 3 0 3 0 2 3 1 0
2 3 3
8 3 3 0 2 1 2 0 0
7 3 1 3 1 3 3 3
11 3 0 3 1 2 0 1 1 3 0 0
3 3 1 3
8 3 0 3 1 3 1 1 1
1 3
12 3 3 2 0 1 1 1 2 0 2 3 1
19 3 1 1 3 3 0 0 3 1 2 1 1 1 2 3 0 1 3 3
6 3 0 2 3 1 2
8 3 3 0 0 1 1 3 0
6 3 2 0 3 1 3
2 3 3
6 3 0 3 0 2 3
3 3 1 3
22 3 1 3 0 2 0 3 1 0 1 3 3 3 1 3 3 0 3 1 2 2 0
4 3 3 2 3
1 3
2 3 3
3 3 3 2
10 3 3 1 3 3 1 3 0 0 0
4 3 3 0 3
9 3 0 3 1 0 1 2 1 3
9 3 3 1 3 0 3 1 3 3
2 3 1
3 3 3 0
2 3 3
5 3 0 3 0 2
18 3 0 3 1 3 3 1 3 3 3 1 0 2 3 1 2 0 0
7 3 3 1 2 1 1 1
3 3 0 3
4 3 0 2 3
22 3 0 3 0 0 2 3 0 3 1 2 1 1 1 3 3 3 3 1 3 0 0
10 3 0 3 0 2 1 0 1 2 3
2 3 0
5 3 3 1 0 0
1 3
6 3 0 3 0 0 2
19 3 1 1 1 1 3 3 0 1 2 3 0 2 1 1 1 1 1 1
2 3 3
10 3 0 3 1 3 3 1 3 0 3
2 3 3
5 3 1 1 3 3
30 3 1 1 1 3 0 2 0 3 1 0 1 2 3 0 3 1 2 1 2 0 2 0 1 0 0 2 0 2 3
9 3 0 3 0 1 3 0 2 3
16 3 0 3 1 3 0 2 3 0 2 0 3 0 1 3 3
15 3 3 0 3 3 1 0 1 3 3 1 3 1 3 3
12 3 3 3 1 3 0 3 0 3 0 3 3
7 3 0 3 1 1 3 0
16 3 0 3 1 2 3 0 1 1 2 1 3 2 1 3 0
14 3 0 3 0 3 1 2 0 3 0 1 1 0 2
22 3 0 3 0 1 0 1 2 3 1 3 0 1 1 1 0 1 3 3 3 3 0
4 3 3 0 0
4 3 1 1 3
13 3 3 0 2 0 3 1 2 1 2 0 2 0
24 3 0 3 0 2 3 0 1 1 1 2 0 3 1 2 1 1 1 2 0 3 2 0 3
1 3
7 3 0 3 0 1 0 2
7 3 0 2 1 1 1 3
2 3 0
9 3 0 2 0 1 3 3 0 2
3 3 3 2
5 3 3 1 3 3
7 3 1 3 0 2 3 3
3 3 0 3
8 3 0 3 0 3 1 2 1
2 3 0
5 3 1 1 3 0
8 3 3 0 3 3 0 3 3
5 3 0 3 3 0
1 3
8 3 0 3 1 2 0 1 3
9 3 0 3 1 0 1 2 0 3
1 3
2 3 3
15 3 3 0 2 0 2 3 1 2 3 1 3 0 0 0
3 3 3 0
10 3 3 0 2 3 1 2 3 3 0
15 3 0 3 1 0 1 3 3 0 3 1 3 0 1 3
7 3 0 2 1 3 0 2
1 3
3 3 3 0
6 3 0 3 1 2 1
21 3 0 3 0 1 3 3 1 3 0 3 1 0 2 1 1 0 0 0 3 1
15 3 0 3 0 2 1 3 0 0 2 0 3 1 0 2
4 3 3 1 2
12 3 0 3 1 3 0 3 0 3 0 2 0
4 3 0 3 0
16 3 0 3 1 3 3 1 1 3 0 0 2 3 0 1 1
7 3 1 3 0 2 3 0
4 3 3 3 3
2 3 3
2 3 0
7 3 1 3 2 3 1 0
2 3 3
3 3 1 3