2566 47
13 1 2 2 2 2 3 4 5 6 7 8 9 10 
11 1 4 5 6 11 12 13 14 15 16 17 
12 1 4 5 6 11 12 13 14 18 19 20 21 
20 1 4 5 6 11 12 13 14 11 12 13 14 22 23 24 25 7 8 9 10 
20 1 4 5 6 11 12 13 14 11 12 13 14 22 23 26 24 25 15 16 17 
19 1 4 5 6 11 12 13 14 11 12 13 14 22 23 24 25 15 16 17 
19 1 4 5 6 11 12 13 14 11 12 13 14 22 23 26 24 25 27 28 
18 1 4 5 6 11 12 13 14 11 12 13 14 22 23 24 25 27 28 
17 1 4 5 6 11 12 13 14 11 12 13 14 15 16 17 8 10 
18 1 4 5 6 11 12 13 14 11 12 13 14 15 16 17 15 16 17 
19 1 4 5 6 11 12 13 14 11 12 13 14 15 16 17 7 27 9 28 
20 1 4 5 6 11 12 13 14 11 12 13 14 15 16 17 29 7 20 9 21 
18 1 4 5 6 11 12 13 14 11 12 13 14 27 28 7 8 9 10 
14 1 4 5 6 11 12 13 14 30 31 7 8 9 10 
17 1 4 5 6 11 12 13 14 11 12 13 14 27 28 15 16 17 
16 1 4 5 6 11 12 13 14 11 12 13 14 27 28 27 28 
18 1 4 5 6 11 12 13 14 11 12 13 14 13 32 7 8 9 10 
17 1 4 5 6 11 12 13 14 11 12 13 14 13 32 15 16 17 
16 1 4 5 6 11 12 13 14 11 12 13 14 13 32 27 28 
17 1 4 5 6 11 12 13 14 11 12 13 14 33 7 8 9 10 
15 1 4 5 6 11 12 13 14 11 12 13 14 33 27 28 
18 1 4 5 6 11 12 13 14 11 12 13 14 34 35 7 8 9 10 
17 1 4 5 6 11 12 13 14 11 12 13 14 34 35 15 16 17 
16 1 4 5 6 11 12 13 14 11 12 13 14 34 35 27 28 
13 1 4 5 6 11 12 13 14 30 31 15 16 17 
16 1 4 5 6 11 12 13 14 11 12 13 14 34 35 20 21 
18 1 4 5 6 11 12 13 14 11 12 13 14 36 37 7 8 9 10 
17 1 4 5 6 11 12 13 14 11 12 13 14 36 37 15 16 17 
16 1 4 5 6 11 12 13 14 11 12 13 14 36 37 27 28 
16 1 4 5 6 11 12 13 14 11 12 13 14 36 37 20 21 
18 1 4 5 6 11 12 13 14 11 12 13 14 38 39 7 8 9 10 
17 1 4 5 6 11 12 13 14 11 12 13 14 38 39 15 16 17 
16 1 4 5 6 11 12 13 14 11 12 13 14 38 39 27 28 
17 1 4 5 6 11 12 13 14 11 12 13 14 40 7 8 9 10 
15 1 4 5 6 11 12 13 14 11 12 13 14 40 27 28 
12 1 4 5 6 11 12 13 14 30 31 27 28 
18 1 4 5 6 11 12 13 14 11 12 13 14 20 21 7 8 9 10 
17 1 4 5 6 11 12 13 14 11 12 13 14 20 21 15 16 17 
16 1 4 5 6 11 12 13 14 11 12 13 14 20 21 27 28 
16 1 4 5 6 11 12 13 14 11 12 13 14 20 21 20 21 
15 1 4 5 6 11 12 13 14 41 42 43 7 8 9 10 
13 1 4 5 6 11 12 13 14 41 42 43 27 28 
14 1 4 5 6 11 12 13 14 41 41 7 8 9 10 
13 1 4 5 6 11 12 13 14 41 41 15 16 17 
12 1 4 5 6 11 12 13 14 41 41 27 28 
15 1 4 5 6 11 12 13 14 41 44 45 7 8 9 10 
12 1 4 5 6 11 12 13 14 30 31 20 21 
13 1 4 5 6 11 12 13 14 41 44 45 27 28 
15 1 4 5 6 11 12 13 14 41 30 31 7 8 9 10 
14 1 4 5 6 11 12 13 14 41 30 31 15 16 17 
13 1 4 5 6 11 12 13 14 41 30 31 27 28 
13 1 4 5 6 11 12 13 14 41 30 31 20 21 
15 1 4 5 6 11 12 13 14 41 46 47 7 8 9 10 
13 1 4 5 6 11 12 13 14 41 46 47 27 28 
13 1 4 5 6 11 12 13 14 41 46 47 20 21 
14 1 4 5 6 11 12 13 14 41 15 16 17 8 10 
15 1 4 5 6 11 12 13 14 41 15 16 17 15 16 17 
14 1 4 5 6 11 12 13 14 46 47 7 8 9 10 
16 1 4 5 6 11 12 13 14 41 15 16 17 7 27 9 28 
17 1 4 5 6 11 12 13 14 41 15 16 17 29 7 20 9 21 
15 1 4 5 6 11 12 13 14 41 27 28 7 8 9 10 
14 1 4 5 6 11 12 13 14 41 27 28 15 16 17 
13 1 4 5 6 11 12 13 14 41 27 28 27 28 
14 1 4 5 6 11 12 13 14 41 33 7 8 9 10 
12 1 4 5 6 11 12 13 14 41 33 27 28 
15 1 4 5 6 11 12 13 14 41 38 39 7 8 9 10 
14 1 4 5 6 11 12 13 14 41 38 39 15 16 17 
13 1 4 5 6 11 12 13 14 41 38 39 27 28 
13 1 4 5 6 11 12 13 14 46 47 15 16 17 
14 1 4 5 6 11 12 13 14 41 40 7 8 9 10 
12 1 4 5 6 11 12 13 14 41 40 27 28 
16 1 4 5 6 11 12 13 14 44 45 42 43 7 8 9 10 
14 1 4 5 6 11 12 13 14 44 45 42 43 27 28 
18 1 4 5 6 11 12 13 14 44 45 11 12 13 14 7 8 9 10 
17 1 4 5 6 11 12 13 14 44 45 11 12 13 14 15 16 17 
16 1 4 5 6 11 12 13 14 44 45 11 12 13 14 27 28 
16 1 4 5 6 11 12 13 14 44 45 11 12 13 14 20 21 
16 1 4 5 6 11 12 13 14 44 45 44 45 7 8 9 10 
14 1 4 5 6 11 12 13 14 44 45 44 45 27 28 
12 1 4 5 6 11 12 13 14 46 47 27 28 
19 1 4 5 6 11 12 13 14 44 45 22 23 26 24 25 7 8 9 10 
18 1 4 5 6 11 12 13 14 44 45 22 23 24 25 7 8 9 10 
18 1 4 5 6 11 12 13 14 44 45 22 23 26 24 25 15 16 17 
17 1 4 5 6 11 12 13 14 44 45 22 23 24 25 15 16 17 
17 1 4 5 6 11 12 13 14 44 45 22 23 26 24 25 27 28 
16 1 4 5 6 11 12 13 14 44 45 22 23 24 25 27 28 
16 1 4 5 6 11 12 13 14 44 45 27 28 7 8 9 10 
15 1 4 5 6 11 12 13 14 44 45 27 28 15 16 17 
14 1 4 5 6 11 12 13 14 44 45 27 28 27 28 
16 1 4 5 6 11 12 13 14 44 45 34 35 7 8 9 10 
12 1 4 5 6 11 12 13 14 46 47 20 21 
15 1 4 5 6 11 12 13 14 44 45 34 35 15 16 17 
14 1 4 5 6 11 12 13 14 44 45 34 35 27 28 
14 1 4 5 6 11 12 13 14 44 45 34 35 20 21 
16 1 4 5 6 11 12 13 14 18 19 42 43 7 8 9 10 
14 1 4 5 6 11 12 13 14 18 19 42 43 27 28 
15 1 4 5 6 11 12 13 14 18 19 41 7 8 9 10 
14 1 4 5 6 11 12 13 14 18 19 41 15 16 17 
13 1 4 5 6 11 12 13 14 18 19 41 27 28 
16 1 4 5 6 11 12 13 14 18 19 44 45 7 8 9 10 
14 1 4 5 6 11 12 13 14 18 19 44 45 27 28 
17 1 4 5 6 11 12 13 14 22 23 26 24 25 7 8 9 10 
16 1 4 5 6 11 12 13 14 18 19 18 19 7 8 9 10 
15 1 4 5 6 11 12 13 14 18 19 18 19 15 16 17 
14 1 4 5 6 11 12 13 14 18 19 18 19 27 28 
14 1 4 5 6 11 12 13 14 18 19 18 19 20 21 
16 1 4 5 6 11 12 13 14 18 19 30 31 7 8 9 10 
15 1 4 5 6 11 12 13 14 18 19 30 31 15 16 17 
14 1 4 5 6 11 12 13 14 18 19 30 31 27 28 
14 1 4 5 6 11 12 13 14 18 19 30 31 20 21 
16 1 4 5 6 11 12 13 14 18 19 46 47 7 8 9 10 
14 1 4 5 6 11 12 13 14 18 19 46 47 27 28 
10 1 4 5 6 11 12 13 14 27 28 
16 1 4 5 6 11 12 13 14 22 23 24 25 7 8 9 10 
14 1 4 5 6 11 12 13 14 18 19 46 47 20 21 
19 1 4 5 6 11 12 13 14 18 19 22 23 26 24 25 7 8 9 10 
18 1 4 5 6 11 12 13 14 18 19 22 23 24 25 7 8 9 10 
18 1 4 5 6 11 12 13 14 18 19 22 23 26 24 25 15 16 17 
17 1 4 5 6 11 12 13 14 18 19 22 23 24 25 15 16 17 
17 1 4 5 6 11 12 13 14 18 19 22 23 26 24 25 27 28 
16 1 4 5 6 11 12 13 14 18 19 22 23 24 25 27 28 
15 1 4 5 6 11 12 13 14 18 19 15 16 17 8 10 
16 1 4 5 6 11 12 13 14 18 19 15 16 17 15 16 17 
17 1 4 5 6 11 12 13 14 18 19 15 16 17 7 27 9 28 
16 1 4 5 6 11 12 13 14 22 23 26 24 25 15 16 17 
18 1 4 5 6 11 12 13 14 18 19 15 16 17 29 7 20 9 21 
16 1 4 5 6 11 12 13 14 18 19 27 28 7 8 9 10 
15 1 4 5 6 11 12 13 14 18 19 27 28 15 16 17 
14 1 4 5 6 11 12 13 14 18 19 27 28 27 28 
16 1 4 5 6 11 12 13 14 18 19 13 32 7 8 9 10 
15 1 4 5 6 11 12 13 14 18 19 13 32 15 16 17 
14 1 4 5 6 11 12 13 14 18 19 13 32 27 28 
15 1 4 5 6 11 12 13 14 18 19 33 7 8 9 10 
13 1 4 5 6 11 12 13 14 18 19 33 27 28 
16 1 4 5 6 11 12 13 14 18 19 36 37 7 8 9 10 
15 1 4 5 6 11 12 13 14 22 23 24 25 15 16 17 
15 1 4 5 6 11 12 13 14 18 19 36 37 15 16 17 
14 1 4 5 6 11 12 13 14 18 19 36 37 27 28 
14 1 4 5 6 11 12 13 14 18 19 36 37 20 21 
16 1 4 5 6 11 12 13 14 18 19 38 39 7 8 9 10 
15 1 4 5 6 11 12 13 14 18 19 38 39 15 16 17 
14 1 4 5 6 11 12 13 14 18 19 38 39 27 28 
15 1 4 5 6 11 12 13 14 18 19 40 7 8 9 10 
13 1 4 5 6 11 12 13 14 18 19 40 27 28 
16 1 4 5 6 11 12 13 14 18 19 20 21 7 8 9 10 
15 1 4 5 6 11 12 13 14 18 19 20 21 15 16 17 
15 1 4 5 6 11 12 13 14 22 23 26 24 25 27 28 
14 1 4 5 6 11 12 13 14 18 19 20 21 27 28 
14 1 4 5 6 11 12 13 14 18 19 20 21 20 21 
16 1 4 5 6 11 12 13 14 30 31 42 43 7 8 9 10 
14 1 4 5 6 11 12 13 14 30 31 42 43 27 28 
16 1 4 5 6 11 12 13 14 30 31 44 45 7 8 9 10 
14 1 4 5 6 11 12 13 14 30 31 44 45 27 28 
16 1 4 5 6 11 12 13 14 30 31 30 31 7 8 9 10 
15 1 4 5 6 11 12 13 14 30 31 30 31 15 16 17 
14 1 4 5 6 11 12 13 14 30 31 30 31 27 28 
14 1 4 5 6 11 12 13 14 30 31 30 31 20 21 
14 1 4 5 6 11 12 13 14 22 23 24 25 27 28 
16 1 4 5 6 11 12 13 14 30 31 46 47 7 8 9 10 
14 1 4 5 6 11 12 13 14 30 31 46 47 27 28 
14 1 4 5 6 11 12 13 14 30 31 46 47 20 21 
19 1 4 5 6 11 12 13 14 30 31 22 23 26 24 25 7 8 9 10 
18 1 4 5 6 11 12 13 14 30 31 22 23 24 25 7 8 9 10 
18 1 4 5 6 11 12 13 14 30 31 22 23 26 24 25 15 16 17 
17 1 4 5 6 11 12 13 14 30 31 22 23 24 25 15 16 17 
17 1 4 5 6 11 12 13 14 30 31 22 23 26 24 25 27 28 
16 1 4 5 6 11 12 13 14 30 31 22 23 24 25 27 28 
15 1 4 5 6 11 12 13 14 30 31 15 16 17 8 10 
15 1 4 5 6 11 12 13 14 22 23 26 24 25 20 21 
16 1 4 5 6 11 12 13 14 30 31 15 16 17 15 16 17 
17 1 4 5 6 11 12 13 14 30 31 15 16 17 7 27 9 28 
18 1 4 5 6 11 12 13 14 30 31 15 16 17 29 7 20 9 21 
16 1 4 5 6 11 12 13 14 30 31 27 28 7 8 9 10 
15 1 4 5 6 11 12 13 14 30 31 27 28 15 16 17 
14 1 4 5 6 11 12 13 14 30 31 27 28 27 28 
15 1 4 5 6 11 12 13 14 30 31 33 7 8 9 10 
13 1 4 5 6 11 12 13 14 30 31 33 27 28 
15 1 4 5 6 11 12 13 14 30 31 40 7 8 9 10 
13 1 4 5 6 11 12 13 14 30 31 40 27 28 
14 1 4 5 6 11 12 13 14 22 23 24 25 20 21 
16 1 4 5 6 11 12 13 14 30 31 20 21 7 8 9 10 
15 1 4 5 6 11 12 13 14 30 31 20 21 15 16 17 
14 1 4 5 6 11 12 13 14 30 31 20 21 27 28 
14 1 4 5 6 11 12 13 14 30 31 20 21 20 21 
16 1 4 5 6 11 12 13 14 46 47 42 43 7 8 9 10 
14 1 4 5 6 11 12 13 14 46 47 42 43 27 28 
18 1 4 5 6 11 12 13 14 46 47 11 12 13 14 7 8 9 10 
17 1 4 5 6 11 12 13 14 46 47 11 12 13 14 15 16 17 
16 1 4 5 6 11 12 13 14 46 47 11 12 13 14 27 28 
16 1 4 5 6 11 12 13 14 46 47 11 12 13 14 20 21 
13 1 4 5 6 11 12 13 14 15 16 17 8 10 
16 1 4 5 6 11 12 13 14 46 47 44 45 7 8 9 10 
14 1 4 5 6 11 12 13 14 46 47 44 45 27 28 
16 1 4 5 6 11 12 13 14 46 47 46 47 7 8 9 10 
14 1 4 5 6 11 12 13 14 46 47 46 47 27 28 
14 1 4 5 6 11 12 13 14 46 47 46 47 20 21 
19 1 4 5 6 11 12 13 14 46 47 22 23 26 24 25 7 8 9 10 
18 1 4 5 6 11 12 13 14 46 47 22 23 24 25 7 8 9 10 
18 1 4 5 6 11 12 13 14 46 47 22 23 26 24 25 15 16 17 
17 1 4 5 6 11 12 13 14 46 47 22 23 24 25 15 16 17 
17 1 4 5 6 11 12 13 14 46 47 22 23 26 24 25 27 28 
14 1 4 5 6 11 12 13 14 15 16 17 15 16 17 
16 1 4 5 6 11 12 13 14 46 47 22 23 24 25 27 28 
16 1 4 5 6 11 12 13 14 46 47 27 28 7 8 9 10 
15 1 4 5 6 11 12 13 14 46 47 27 28 15 16 17 
14 1 4 5 6 11 12 13 14 46 47 27 28 27 28 
16 1 4 5 6 11 12 13 14 46 47 34 35 7 8 9 10 
15 1 4 5 6 11 12 13 14 46 47 34 35 15 16 17 
14 1 4 5 6 11 12 13 14 46 47 34 35 27 28 
14 1 4 5 6 11 12 13 14 46 47 34 35 20 21 
15 1 4 5 6 11 12 13 14 46 47 40 7 8 9 10 
13 1 4 5 6 11 12 13 14 46 47 40 27 28 
15 1 4 5 6 11 12 13 14 15 16 17 7 27 9 28 
16 1 4 5 6 11 12 13 14 46 47 20 21 7 8 9 10 
15 1 4 5 6 11 12 13 14 46 47 20 21 15 16 17 
14 1 4 5 6 11 12 13 14 46 47 20 21 27 28 
14 1 4 5 6 11 12 13 14 46 47 20 21 20 21 
19 1 4 5 6 11 12 13 14 22 23 26 24 25 42 43 7 8 9 10 
18 1 4 5 6 11 12 13 14 22 23 24 25 42 43 7 8 9 10 
17 1 4 5 6 11 12 13 14 22 23 26 24 25 42 43 27 28 
16 1 4 5 6 11 12 13 14 22 23 24 25 42 43 27 28 
21 1 4 5 6 11 12 13 14 22 23 26 24 25 11 12 13 14 7 8 9 10 
20 1 4 5 6 11 12 13 14 22 23 24 25 11 12 13 14 7 8 9 10 
10 1 4 5 6 11 12 13 14 20 21 
16 1 4 5 6 11 12 13 14 15 16 17 29 7 20 9 21 
20 1 4 5 6 11 12 13 14 22 23 26 24 25 11 12 13 14 15 16 17 
19 1 4 5 6 11 12 13 14 22 23 24 25 11 12 13 14 15 16 17 
19 1 4 5 6 11 12 13 14 22 23 26 24 25 11 12 13 14 27 28 
18 1 4 5 6 11 12 13 14 22 23 24 25 11 12 13 14 27 28 
19 1 4 5 6 11 12 13 14 22 23 26 24 25 11 12 13 14 20 21 
18 1 4 5 6 11 12 13 14 22 23 24 25 11 12 13 14 20 21 
18 1 4 5 6 11 12 13 14 22 23 26 24 25 41 7 8 9 10 
17 1 4 5 6 11 12 13 14 22 23 24 25 41 7 8 9 10 
17 1 4 5 6 11 12 13 14 22 23 26 24 25 41 15 16 17 
16 1 4 5 6 11 12 13 14 22 23 24 25 41 15 16 17 
14 1 4 5 6 11 12 13 14 27 28 7 8 9 10 
16 1 4 5 6 11 12 13 14 22 23 26 24 25 41 27 28 
15 1 4 5 6 11 12 13 14 22 23 24 25 41 27 28 
19 1 4 5 6 11 12 13 14 22 23 26 24 25 44 45 7 8 9 10 
18 1 4 5 6 11 12 13 14 22 23 24 25 44 45 7 8 9 10 
17 1 4 5 6 11 12 13 14 22 23 26 24 25 44 45 27 28 
16 1 4 5 6 11 12 13 14 22 23 24 25 44 45 27 28 
19 1 4 5 6 11 12 13 14 22 23 26 24 25 18 19 7 8 9 10 
18 1 4 5 6 11 12 13 14 22 23 24 25 18 19 7 8 9 10 
18 1 4 5 6 11 12 13 14 22 23 26 24 25 18 19 15 16 17 
17 1 4 5 6 11 12 13 14 22 23 24 25 18 19 15 16 17 
13 1 4 5 6 11 12 13 14 27 28 15 16 17 
17 1 4 5 6 11 12 13 14 22 23 26 24 25 18 19 27 28 
16 1 4 5 6 11 12 13 14 22 23 24 25 18 19 27 28 
17 1 4 5 6 11 12 13 14 22 23 26 24 25 18 19 20 21 
16 1 4 5 6 11 12 13 14 22 23 24 25 18 19 20 21 
19 1 4 5 6 11 12 13 14 22 23 26 24 25 30 31 7 8 9 10 
18 1 4 5 6 11 12 13 14 22 23 24 25 30 31 7 8 9 10 
18 1 4 5 6 11 12 13 14 22 23 26 24 25 30 31 15 16 17 
17 1 4 5 6 11 12 13 14 22 23 24 25 30 31 15 16 17 
17 1 4 5 6 11 12 13 14 22 23 26 24 25 30 31 27 28 
16 1 4 5 6 11 12 13 14 22 23 24 25 30 31 27 28 
12 1 4 5 6 11 12 13 14 27 28 27 28 
17 1 4 5 6 11 12 13 14 22 23 26 24 25 30 31 20 21 
16 1 4 5 6 11 12 13 14 22 23 24 25 30 31 20 21 
19 1 4 5 6 11 12 13 14 22 23 26 24 25 46 47 7 8 9 10 
18 1 4 5 6 11 12 13 14 22 23 24 25 46 47 7 8 9 10 
17 1 4 5 6 11 12 13 14 22 23 26 24 25 46 47 27 28 
16 1 4 5 6 11 12 13 14 22 23 24 25 46 47 27 28 
17 1 4 5 6 11 12 13 14 22 23 26 24 25 46 47 20 21 
16 1 4 5 6 11 12 13 14 22 23 24 25 46 47 20 21 
22 1 4 5 6 11 12 13 14 22 23 26 24 25 22 23 26 24 25 7 8 9 10 
21 1 4 5 6 11 12 13 14 22 23 26 24 25 22 23 24 25 7 8 9 10 
12 1 4 5 6 11 12 13 14 27 28 20 21 
21 1 4 5 6 11 12 13 14 22 23 24 25 22 23 26 24 25 7 8 9 10 
20 1 4 5 6 11 12 13 14 22 23 24 25 22 23 24 25 7 8 9 10 
21 1 4 5 6 11 12 13 14 22 23 26 24 25 22 23 26 24 25 15 16 17 
20 1 4 5 6 11 12 13 14 22 23 26 24 25 22 23 24 25 15 16 17 
20 1 4 5 6 11 12 13 14 22 23 24 25 22 23 26 24 25 15 16 17 
19 1 4 5 6 11 12 13 14 22 23 24 25 22 23 24 25 15 16 17 
20 1 4 5 6 11 12 13 14 22 23 26 24 25 22 23 26 24 25 27 28 
19 1 4 5 6 11 12 13 14 22 23 26 24 25 22 23 24 25 27 28 
19 1 4 5 6 11 12 13 14 22 23 24 25 22 23 26 24 25 27 28 
18 1 4 5 6 11 12 13 14 22 23 24 25 22 23 24 25 27 28 
14 1 4 5 6 11 12 13 14 13 32 7 8 9 10 
18 1 4 5 6 11 12 13 14 22 23 26 24 25 15 16 17 8 10 
17 1 4 5 6 11 12 13 14 22 23 24 25 15 16 17 8 10 
19 1 4 5 6 11 12 13 14 22 23 26 24 25 15 16 17 15 16 17 
18 1 4 5 6 11 12 13 14 22 23 24 25 15 16 17 15 16 17 
20 1 4 5 6 11 12 13 14 22 23 26 24 25 15 16 17 7 27 9 28 
19 1 4 5 6 11 12 13 14 22 23 24 25 15 16 17 7 27 9 28 
21 1 4 5 6 11 12 13 14 22 23 26 24 25 15 16 17 29 7 20 9 21 
20 1 4 5 6 11 12 13 14 22 23 24 25 15 16 17 29 7 20 9 21 
19 1 4 5 6 11 12 13 14 22 23 26 24 25 27 28 7 8 9 10 
18 1 4 5 6 11 12 13 14 22 23 24 25 27 28 7 8 9 10 
13 1 4 5 6 11 12 13 14 13 32 15 16 17 
18 1 4 5 6 11 12 13 14 22 23 26 24 25 27 28 15 16 17 
17 1 4 5 6 11 12 13 14 22 23 24 25 27 28 15 16 17 
17 1 4 5 6 11 12 13 14 22 23 26 24 25 27 28 27 28 
16 1 4 5 6 11 12 13 14 22 23 24 25 27 28 27 28 
19 1 4 5 6 11 12 13 14 22 23 26 24 25 13 32 7 8 9 10 
18 1 4 5 6 11 12 13 14 22 23 24 25 13 32 7 8 9 10 
18 1 4 5 6 11 12 13 14 22 23 26 24 25 13 32 15 16 17 
17 1 4 5 6 11 12 13 14 22 23 24 25 13 32 15 16 17 
17 1 4 5 6 11 12 13 14 22 23 26 24 25 13 32 27 28 
16 1 4 5 6 11 12 13 14 22 23 24 25 13 32 27 28 
12 1 4 5 6 11 12 13 14 13 32 27 28 
18 1 4 5 6 11 12 13 14 22 23 26 24 25 33 7 8 9 10 
17 1 4 5 6 11 12 13 14 22 23 24 25 33 7 8 9 10 
16 1 4 5 6 11 12 13 14 22 23 26 24 25 33 27 28 
15 1 4 5 6 11 12 13 14 22 23 24 25 33 27 28 
19 1 4 5 6 11 12 13 14 22 23 26 24 25 34 35 7 8 9 10 
18 1 4 5 6 11 12 13 14 22 23 24 25 34 35 7 8 9 10 
18 1 4 5 6 11 12 13 14 22 23 26 24 25 34 35 15 16 17 
17 1 4 5 6 11 12 13 14 22 23 24 25 34 35 15 16 17 
17 1 4 5 6 11 12 13 14 22 23 26 24 25 34 35 27 28 
16 1 4 5 6 11 12 13 14 22 23 24 25 34 35 27 28 
12 1 4 5 6 11 12 13 14 13 32 20 21 
17 1 4 5 6 11 12 13 14 22 23 26 24 25 34 35 20 21 
16 1 4 5 6 11 12 13 14 22 23 24 25 34 35 20 21 
19 1 4 5 6 11 12 13 14 22 23 26 24 25 36 37 7 8 9 10 
18 1 4 5 6 11 12 13 14 22 23 24 25 36 37 7 8 9 10 
18 1 4 5 6 11 12 13 14 22 23 26 24 25 36 37 15 16 17 
17 1 4 5 6 11 12 13 14 22 23 24 25 36 37 15 16 17 
17 1 4 5 6 11 12 13 14 22 23 26 24 25 36 37 27 28 
16 1 4 5 6 11 12 13 14 22 23 24 25 36 37 27 28 
17 1 4 5 6 11 12 13 14 22 23 26 24 25 36 37 20 21 
16 1 4 5 6 11 12 13 14 22 23 24 25 36 37 20 21 
13 1 4 5 6 11 12 13 14 33 7 8 9 10 
19 1 4 5 6 11 12 13 14 22 23 26 24 25 38 39 7 8 9 10 
18 1 4 5 6 11 12 13 14 22 23 24 25 38 39 7 8 9 10 
18 1 4 5 6 11 12 13 14 22 23 26 24 25 38 39 15 16 17 
17 1 4 5 6 11 12 13 14 22 23 24 25 38 39 15 16 17 
17 1 4 5 6 11 12 13 14 22 23 26 24 25 38 39 27 28 
16 1 4 5 6 11 12 13 14 22 23 24 25 38 39 27 28 
18 1 4 5 6 11 12 13 14 22 23 26 24 25 40 7 8 9 10 
17 1 4 5 6 11 12 13 14 22 23 24 25 40 7 8 9 10 
16 1 4 5 6 11 12 13 14 22 23 26 24 25 40 27 28 
15 1 4 5 6 11 12 13 14 22 23 24 25 40 27 28 
8 1 4 5 6 7 8 9 10 
12 1 4 5 6 11 12 13 14 33 15 16 17 
16 1 4 5 6 11 12 13 14 27 28 30 31 7 8 9 10 
15 1 4 5 6 11 12 13 14 27 28 30 31 15 16 17 
14 1 4 5 6 11 12 13 14 27 28 30 31 27 28 
14 1 4 5 6 11 12 13 14 27 28 30 31 20 21 
15 1 4 5 6 11 12 13 14 27 28 15 16 17 8 10 
16 1 4 5 6 11 12 13 14 27 28 15 16 17 15 16 17 
17 1 4 5 6 11 12 13 14 27 28 15 16 17 7 27 9 28 
18 1 4 5 6 11 12 13 14 27 28 15 16 17 29 7 20 9 21 
16 1 4 5 6 11 12 13 14 27 28 27 28 7 8 9 10 
15 1 4 5 6 11 12 13 14 27 28 27 28 15 16 17 
11 1 4 5 6 11 12 13 14 33 27 28 
14 1 4 5 6 11 12 13 14 27 28 27 28 27 28 
16 1 4 5 6 11 12 13 14 27 28 38 39 7 8 9 10 
15 1 4 5 6 11 12 13 14 27 28 38 39 15 16 17 
14 1 4 5 6 11 12 13 14 27 28 38 39 27 28 
16 1 4 5 6 11 12 13 14 13 32 42 43 7 8 9 10 
14 1 4 5 6 11 12 13 14 13 32 42 43 27 28 
15 1 4 5 6 11 12 13 14 13 32 41 7 8 9 10 
14 1 4 5 6 11 12 13 14 13 32 41 15 16 17 
13 1 4 5 6 11 12 13 14 13 32 41 27 28 
16 1 4 5 6 11 12 13 14 13 32 44 45 7 8 9 10 
11 1 4 5 6 11 12 13 14 33 20 21 
14 1 4 5 6 11 12 13 14 13 32 44 45 27 28 
16 1 4 5 6 11 12 13 14 13 32 30 31 7 8 9 10 
15 1 4 5 6 11 12 13 14 13 32 30 31 15 16 17 
14 1 4 5 6 11 12 13 14 13 32 30 31 27 28 
14 1 4 5 6 11 12 13 14 13 32 30 31 20 21 
16 1 4 5 6 11 12 13 14 13 32 46 47 7 8 9 10 
14 1 4 5 6 11 12 13 14 13 32 46 47 27 28 
14 1 4 5 6 11 12 13 14 13 32 46 47 20 21 
15 1 4 5 6 11 12 13 14 13 32 15 16 17 8 10 
16 1 4 5 6 11 12 13 14 13 32 15 16 17 15 16 17 
14 1 4 5 6 11 12 13 14 34 35 7 8 9 10 
17 1 4 5 6 11 12 13 14 13 32 15 16 17 7 27 9 28 
18 1 4 5 6 11 12 13 14 13 32 15 16 17 29 7 20 9 21 
16 1 4 5 6 11 12 13 14 13 32 27 28 7 8 9 10 
15 1 4 5 6 11 12 13 14 13 32 27 28 15 16 17 
14 1 4 5 6 11 12 13 14 13 32 27 28 27 28 
16 1 4 5 6 11 12 13 14 13 32 13 32 7 8 9 10 
15 1 4 5 6 11 12 13 14 13 32 13 32 15 16 17 
14 1 4 5 6 11 12 13 14 13 32 13 32 27 28 
15 1 4 5 6 11 12 13 14 13 32 33 7 8 9 10 
13 1 4 5 6 11 12 13 14 13 32 33 27 28 
13 1 4 5 6 11 12 13 14 34 35 15 16 17 
16 1 4 5 6 11 12 13 14 13 32 36 37 7 8 9 10 
15 1 4 5 6 11 12 13 14 13 32 36 37 15 16 17 
14 1 4 5 6 11 12 13 14 13 32 36 37 27 28 
14 1 4 5 6 11 12 13 14 13 32 36 37 20 21 
16 1 4 5 6 11 12 13 14 13 32 38 39 7 8 9 10 
15 1 4 5 6 11 12 13 14 13 32 38 39 15 16 17 
14 1 4 5 6 11 12 13 14 13 32 38 39 27 28 
15 1 4 5 6 11 12 13 14 13 32 40 7 8 9 10 
13 1 4 5 6 11 12 13 14 13 32 40 27 28 
15 1 4 5 6 11 12 13 14 33 42 43 7 8 9 10 
12 1 4 5 6 11 12 13 14 34 35 27 28 
13 1 4 5 6 11 12 13 14 33 42 43 27 28 
15 1 4 5 6 11 12 13 14 33 44 45 7 8 9 10 
13 1 4 5 6 11 12 13 14 33 44 45 27 28 
15 1 4 5 6 11 12 13 14 33 46 47 7 8 9 10 
13 1 4 5 6 11 12 13 14 33 46 47 27 28 
13 1 4 5 6 11 12 13 14 33 46 47 20 21 
15 1 4 5 6 11 12 13 14 33 27 28 7 8 9 10 
14 1 4 5 6 11 12 13 14 33 27 28 15 16 17 
13 1 4 5 6 11 12 13 14 33 27 28 27 28 
14 1 4 5 6 11 12 13 14 33 33 7 8 9 10 
12 1 4 5 6 11 12 13 14 34 35 20 21 
12 1 4 5 6 11 12 13 14 33 33 27 28 
14 1 4 5 6 11 12 13 14 33 40 7 8 9 10 
12 1 4 5 6 11 12 13 14 33 40 27 28 
16 1 4 5 6 11 12 13 14 34 35 42 43 7 8 9 10 
14 1 4 5 6 11 12 13 14 34 35 42 43 27 28 
18 1 4 5 6 11 12 13 14 34 35 11 12 13 14 7 8 9 10 
17 1 4 5 6 11 12 13 14 34 35 11 12 13 14 15 16 17 
16 1 4 5 6 11 12 13 14 34 35 11 12 13 14 27 28 
16 1 4 5 6 11 12 13 14 34 35 11 12 13 14 20 21 
15 1 4 5 6 11 12 13 14 34 35 41 7 8 9 10 
14 1 4 5 6 11 12 13 14 36 37 7 8 9 10 
14 1 4 5 6 11 12 13 14 34 35 41 15 16 17 
13 1 4 5 6 11 12 13 14 34 35 41 27 28 
16 1 4 5 6 11 12 13 14 34 35 44 45 7 8 9 10 
14 1 4 5 6 11 12 13 14 34 35 44 45 27 28 
16 1 4 5 6 11 12 13 14 34 35 18 19 7 8 9 10 
15 1 4 5 6 11 12 13 14 34 35 18 19 15 16 17 
14 1 4 5 6 11 12 13 14 34 35 18 19 27 28 
14 1 4 5 6 11 12 13 14 34 35 18 19 20 21 
16 1 4 5 6 11 12 13 14 34 35 30 31 7 8 9 10 
15 1 4 5 6 11 12 13 14 34 35 30 31 15 16 17 
13 1 4 5 6 11 12 13 14 36 37 15 16 17 
14 1 4 5 6 11 12 13 14 34 35 30 31 27 28 
14 1 4 5 6 11 12 13 14 34 35 30 31 20 21 
16 1 4 5 6 11 12 13 14 34 35 46 47 7 8 9 10 
14 1 4 5 6 11 12 13 14 34 35 46 47 27 28 
14 1 4 5 6 11 12 13 14 34 35 46 47 20 21 
19 1 4 5 6 11 12 13 14 34 35 22 23 26 24 25 7 8 9 10 
18 1 4 5 6 11 12 13 14 34 35 22 23 24 25 7 8 9 10 
18 1 4 5 6 11 12 13 14 34 35 22 23 26 24 25 15 16 17 
17 1 4 5 6 11 12 13 14 34 35 22 23 24 25 15 16 17 
17 1 4 5 6 11 12 13 14 34 35 22 23 26 24 25 27 28 
12 1 4 5 6 11 12 13 14 36 37 27 28 
16 1 4 5 6 11 12 13 14 34 35 22 23 24 25 27 28 
15 1 4 5 6 11 12 13 14 34 35 15 16 17 8 10 
16 1 4 5 6 11 12 13 14 34 35 15 16 17 15 16 17 
17 1 4 5 6 11 12 13 14 34 35 15 16 17 7 27 9 28 
18 1 4 5 6 11 12 13 14 34 35 15 16 17 29 7 20 9 21 
16 1 4 5 6 11 12 13 14 34 35 27 28 7 8 9 10 
15 1 4 5 6 11 12 13 14 34 35 27 28 15 16 17 
14 1 4 5 6 11 12 13 14 34 35 27 28 27 28 
16 1 4 5 6 11 12 13 14 34 35 13 32 7 8 9 10 
15 1 4 5 6 11 12 13 14 34 35 13 32 15 16 17 
8 1 4 5 6 7 8 9 10 
12 1 4 5 6 11 12 13 14 36 37 20 21 
14 1 4 5 6 11 12 13 14 34 35 13 32 27 28 
15 1 4 5 6 11 12 13 14 34 35 33 7 8 9 10 
13 1 4 5 6 11 12 13 14 34 35 33 27 28 
16 1 4 5 6 11 12 13 14 34 35 34 35 7 8 9 10 
15 1 4 5 6 11 12 13 14 34 35 34 35 15 16 17 
14 1 4 5 6 11 12 13 14 34 35 34 35 27 28 
14 1 4 5 6 11 12 13 14 34 35 34 35 20 21 
16 1 4 5 6 11 12 13 14 34 35 36 37 7 8 9 10 
15 1 4 5 6 11 12 13 14 34 35 36 37 15 16 17 
14 1 4 5 6 11 12 13 14 34 35 36 37 27 28 
14 1 4 5 6 11 12 13 14 38 39 7 8 9 10 
14 1 4 5 6 11 12 13 14 34 35 36 37 20 21 
16 1 4 5 6 11 12 13 14 34 35 38 39 7 8 9 10 
15 1 4 5 6 11 12 13 14 34 35 38 39 15 16 17 
14 1 4 5 6 11 12 13 14 34 35 38 39 27 28 
15 1 4 5 6 11 12 13 14 34 35 40 7 8 9 10 
13 1 4 5 6 11 12 13 14 34 35 40 27 28 
16 1 4 5 6 11 12 13 14 34 35 20 21 7 8 9 10 
15 1 4 5 6 11 12 13 14 34 35 20 21 15 16 17 
14 1 4 5 6 11 12 13 14 34 35 20 21 27 28 
14 1 4 5 6 11 12 13 14 34 35 20 21 20 21 
13 1 4 5 6 11 12 13 14 38 39 15 16 17 
16 1 4 5 6 11 12 13 14 36 37 42 43 7 8 9 10 
14 1 4 5 6 11 12 13 14 36 37 42 43 27 28 
18 1 4 5 6 11 12 13 14 36 37 11 12 13 14 7 8 9 10 
17 1 4 5 6 11 12 13 14 36 37 11 12 13 14 15 16 17 
16 1 4 5 6 11 12 13 14 36 37 11 12 13 14 27 28 
16 1 4 5 6 11 12 13 14 36 37 11 12 13 14 20 21 
15 1 4 5 6 11 12 13 14 36 37 41 7 8 9 10 
14 1 4 5 6 11 12 13 14 36 37 41 15 16 17 
13 1 4 5 6 11 12 13 14 36 37 41 27 28 
16 1 4 5 6 11 12 13 14 36 37 44 45 7 8 9 10 
12 1 4 5 6 11 12 13 14 38 39 27 28 
14 1 4 5 6 11 12 13 14 36 37 44 45 27 28 
16 1 4 5 6 11 12 13 14 36 37 30 31 7 8 9 10 
15 1 4 5 6 11 12 13 14 36 37 30 31 15 16 17 
14 1 4 5 6 11 12 13 14 36 37 30 31 27 28 
14 1 4 5 6 11 12 13 14 36 37 30 31 20 21 
16 1 4 5 6 11 12 13 14 36 37 46 47 7 8 9 10 
14 1 4 5 6 11 12 13 14 36 37 46 47 27 28 
14 1 4 5 6 11 12 13 14 36 37 46 47 20 21 
19 1 4 5 6 11 12 13 14 36 37 22 23 26 24 25 7 8 9 10 
18 1 4 5 6 11 12 13 14 36 37 22 23 24 25 7 8 9 10 
12 1 4 5 6 11 12 13 14 38 39 20 21 
18 1 4 5 6 11 12 13 14 36 37 22 23 26 24 25 15 16 17 
17 1 4 5 6 11 12 13 14 36 37 22 23 24 25 15 16 17 
17 1 4 5 6 11 12 13 14 36 37 22 23 26 24 25 27 28 
16 1 4 5 6 11 12 13 14 36 37 22 23 24 25 27 28 
15 1 4 5 6 11 12 13 14 36 37 15 16 17 8 10 
16 1 4 5 6 11 12 13 14 36 37 15 16 17 15 16 17 
17 1 4 5 6 11 12 13 14 36 37 15 16 17 7 27 9 28 
18 1 4 5 6 11 12 13 14 36 37 15 16 17 29 7 20 9 21 
16 1 4 5 6 11 12 13 14 36 37 27 28 7 8 9 10 
15 1 4 5 6 11 12 13 14 36 37 27 28 15 16 17 
13 1 4 5 6 11 12 13 14 40 7 8 9 10 
14 1 4 5 6 11 12 13 14 36 37 27 28 27 28 
15 1 4 5 6 11 12 13 14 36 37 33 7 8 9 10 
13 1 4 5 6 11 12 13 14 36 37 33 27 28 
16 1 4 5 6 11 12 13 14 36 37 34 35 7 8 9 10 
15 1 4 5 6 11 12 13 14 36 37 34 35 15 16 17 
14 1 4 5 6 11 12 13 14 36 37 34 35 27 28 
14 1 4 5 6 11 12 13 14 36 37 34 35 20 21 
16 1 4 5 6 11 12 13 14 36 37 36 37 7 8 9 10 
15 1 4 5 6 11 12 13 14 36 37 36 37 15 16 17 
14 1 4 5 6 11 12 13 14 36 37 36 37 27 28 
12 1 4 5 6 11 12 13 14 40 15 16 17 
14 1 4 5 6 11 12 13 14 36 37 36 37 20 21 
16 1 4 5 6 11 12 13 14 36 37 38 39 7 8 9 10 
15 1 4 5 6 11 12 13 14 36 37 38 39 15 16 17 
14 1 4 5 6 11 12 13 14 36 37 38 39 27 28 
15 1 4 5 6 11 12 13 14 36 37 40 7 8 9 10 
13 1 4 5 6 11 12 13 14 36 37 40 27 28 
16 1 4 5 6 11 12 13 14 36 37 20 21 7 8 9 10 
15 1 4 5 6 11 12 13 14 36 37 20 21 15 16 17 
14 1 4 5 6 11 12 13 14 36 37 20 21 27 28 
14 1 4 5 6 11 12 13 14 36 37 20 21 20 21 
11 1 4 5 6 11 12 13 14 40 27 28 
16 1 4 5 6 11 12 13 14 38 39 42 43 7 8 9 10 
14 1 4 5 6 11 12 13 14 38 39 42 43 27 28 
16 1 4 5 6 11 12 13 14 38 39 44 45 7 8 9 10 
14 1 4 5 6 11 12 13 14 38 39 44 45 27 28 
16 1 4 5 6 11 12 13 14 38 39 30 31 7 8 9 10 
15 1 4 5 6 11 12 13 14 38 39 30 31 15 16 17 
14 1 4 5 6 11 12 13 14 38 39 30 31 27 28 
14 1 4 5 6 11 12 13 14 38 39 30 31 20 21 
16 1 4 5 6 11 12 13 14 38 39 46 47 7 8 9 10 
14 1 4 5 6 11 12 13 14 38 39 46 47 27 28 
11 1 4 5 6 11 12 13 14 40 20 21 
14 1 4 5 6 11 12 13 14 38 39 46 47 20 21 
19 1 4 5 6 11 12 13 14 38 39 22 23 26 24 25 7 8 9 10 
18 1 4 5 6 11 12 13 14 38 39 22 23 24 25 7 8 9 10 
18 1 4 5 6 11 12 13 14 38 39 22 23 26 24 25 15 16 17 
17 1 4 5 6 11 12 13 14 38 39 22 23 24 25 15 16 17 
17 1 4 5 6 11 12 13 14 38 39 22 23 26 24 25 27 28 
16 1 4 5 6 11 12 13 14 38 39 22 23 24 25 27 28 
15 1 4 5 6 11 12 13 14 38 39 15 16 17 8 10 
16 1 4 5 6 11 12 13 14 38 39 15 16 17 15 16 17 
17 1 4 5 6 11 12 13 14 38 39 15 16 17 7 27 9 28 
14 1 4 5 6 11 12 13 14 20 21 7 8 9 10 
18 1 4 5 6 11 12 13 14 38 39 15 16 17 29 7 20 9 21 
16 1 4 5 6 11 12 13 14 38 39 27 28 7 8 9 10 
15 1 4 5 6 11 12 13 14 38 39 27 28 15 16 17 
14 1 4 5 6 11 12 13 14 38 39 27 28 27 28 
15 1 4 5 6 11 12 13 14 38 39 33 7 8 9 10 
13 1 4 5 6 11 12 13 14 38 39 33 27 28 
16 1 4 5 6 11 12 13 14 38 39 38 39 7 8 9 10 
15 1 4 5 6 11 12 13 14 38 39 38 39 15 16 17 
14 1 4 5 6 11 12 13 14 38 39 38 39 27 28 
15 1 4 5 6 11 12 13 14 38 39 40 7 8 9 10 
8 1 4 5 6 7 8 9 10 
13 1 4 5 6 11 12 13 14 20 21 15 16 17 
13 1 4 5 6 11 12 13 14 38 39 40 27 28 
15 1 4 5 6 11 12 13 14 40 42 43 7 8 9 10 
13 1 4 5 6 11 12 13 14 40 42 43 27 28 
15 1 4 5 6 11 12 13 14 40 44 45 7 8 9 10 
13 1 4 5 6 11 12 13 14 40 44 45 27 28 
15 1 4 5 6 11 12 13 14 40 27 28 7 8 9 10 
14 1 4 5 6 11 12 13 14 40 27 28 15 16 17 
13 1 4 5 6 11 12 13 14 40 27 28 27 28 
14 1 4 5 6 11 12 13 14 40 40 7 8 9 10 
12 1 4 5 6 11 12 13 14 40 40 27 28 
12 1 4 5 6 11 12 13 14 20 21 27 28 
16 1 4 5 6 11 12 13 14 20 21 42 43 7 8 9 10 
14 1 4 5 6 11 12 13 14 20 21 42 43 27 28 
18 1 4 5 6 11 12 13 14 20 21 11 12 13 14 7 8 9 10 
17 1 4 5 6 11 12 13 14 20 21 11 12 13 14 15 16 17 
16 1 4 5 6 11 12 13 14 20 21 11 12 13 14 27 28 
16 1 4 5 6 11 12 13 14 20 21 11 12 13 14 20 21 
15 1 4 5 6 11 12 13 14 20 21 41 7 8 9 10 
14 1 4 5 6 11 12 13 14 20 21 41 15 16 17 
13 1 4 5 6 11 12 13 14 20 21 41 27 28 
16 1 4 5 6 11 12 13 14 20 21 44 45 7 8 9 10 
12 1 4 5 6 11 12 13 14 20 21 20 21 
14 1 4 5 6 11 12 13 14 20 21 44 45 27 28 
16 1 4 5 6 11 12 13 14 20 21 18 19 7 8 9 10 
15 1 4 5 6 11 12 13 14 20 21 18 19 15 16 17 
14 1 4 5 6 11 12 13 14 20 21 18 19 27 28 
14 1 4 5 6 11 12 13 14 20 21 18 19 20 21 
16 1 4 5 6 11 12 13 14 20 21 30 31 7 8 9 10 
15 1 4 5 6 11 12 13 14 20 21 30 31 15 16 17 
14 1 4 5 6 11 12 13 14 20 21 30 31 27 28 
14 1 4 5 6 11 12 13 14 20 21 30 31 20 21 
16 1 4 5 6 11 12 13 14 20 21 46 47 7 8 9 10 
12 1 4 5 6 36 37 42 43 7 8 9 10 
14 1 4 5 6 11 12 13 14 20 21 46 47 27 28 
14 1 4 5 6 11 12 13 14 20 21 46 47 20 21 
19 1 4 5 6 11 12 13 14 20 21 22 23 26 24 25 7 8 9 10 
18 1 4 5 6 11 12 13 14 20 21 22 23 24 25 7 8 9 10 
18 1 4 5 6 11 12 13 14 20 21 22 23 26 24 25 15 16 17 
17 1 4 5 6 11 12 13 14 20 21 22 23 24 25 15 16 17 
17 1 4 5 6 11 12 13 14 20 21 22 23 26 24 25 27 28 
16 1 4 5 6 11 12 13 14 20 21 22 23 24 25 27 28 
15 1 4 5 6 11 12 13 14 20 21 15 16 17 8 10 
16 1 4 5 6 11 12 13 14 20 21 15 16 17 15 16 17 
11 1 4 5 6 36 37 42 43 15 16 17 
17 1 4 5 6 11 12 13 14 20 21 15 16 17 7 27 9 28 
18 1 4 5 6 11 12 13 14 20 21 15 16 17 29 7 20 9 21 
16 1 4 5 6 11 12 13 14 20 21 27 28 7 8 9 10 
15 1 4 5 6 11 12 13 14 20 21 27 28 15 16 17 
14 1 4 5 6 11 12 13 14 20 21 27 28 27 28 
16 1 4 5 6 11 12 13 14 20 21 13 32 7 8 9 10 
15 1 4 5 6 11 12 13 14 20 21 13 32 15 16 17 
14 1 4 5 6 11 12 13 14 20 21 13 32 27 28 
15 1 4 5 6 11 12 13 14 20 21 33 7 8 9 10 
13 1 4 5 6 11 12 13 14 20 21 33 27 28 
10 1 4 5 6 36 37 42 43 27 28 
16 1 4 5 6 11 12 13 14 20 21 34 35 7 8 9 10 
15 1 4 5 6 11 12 13 14 20 21 34 35 15 16 17 
14 1 4 5 6 11 12 13 14 20 21 34 35 27 28 
14 1 4 5 6 11 12 13 14 20 21 34 35 20 21 
16 1 4 5 6 11 12 13 14 20 21 36 37 7 8 9 10 
15 1 4 5 6 11 12 13 14 20 21 36 37 15 16 17 
14 1 4 5 6 11 12 13 14 20 21 36 37 27 28 
14 1 4 5 6 11 12 13 14 20 21 36 37 20 21 
16 1 4 5 6 11 12 13 14 20 21 38 39 7 8 9 10 
15 1 4 5 6 11 12 13 14 20 21 38 39 15 16 17 
13 1 4 5 6 36 37 42 43 29 7 20 9 21 
14 1 4 5 6 11 12 13 14 20 21 38 39 27 28 
15 1 4 5 6 11 12 13 14 20 21 40 7 8 9 10 
13 1 4 5 6 11 12 13 14 20 21 40 27 28 
16 1 4 5 6 11 12 13 14 20 21 20 21 7 8 9 10 
15 1 4 5 6 11 12 13 14 20 21 20 21 15 16 17 
14 1 4 5 6 11 12 13 14 20 21 20 21 27 28 
14 1 4 5 6 11 12 13 14 20 21 20 21 20 21 
13 1 4 5 6 41 42 43 42 43 7 8 9 10 
11 1 4 5 6 41 42 43 42 43 27 28 
15 1 4 5 6 41 42 43 11 12 13 14 7 8 9 10 
14 1 4 5 6 36 37 11 12 13 14 7 8 9 10 
14 1 4 5 6 41 42 43 11 12 13 14 15 16 17 
13 1 4 5 6 41 42 43 11 12 13 14 27 28 
13 1 4 5 6 41 42 43 11 12 13 14 20 21 
16 1 4 5 6 41 42 43 22 29 7 23 25 7 8 9 10 
16 1 4 5 6 41 42 43 22 29 7 23 25 7 15 9 17 
14 1 4 5 6 41 42 43 22 29 7 23 25 27 28 
13 1 4 5 6 41 42 43 27 28 7 8 9 10 
13 1 4 5 6 41 42 43 27 28 7 15 9 17 
11 1 4 5 6 41 42 43 27 28 27 28 
13 1 4 5 6 41 42 43 34 35 7 8 9 10 
13 1 4 5 6 36 37 11 12 13 14 15 16 17 
12 1 4 5 6 41 42 43 34 35 15 16 17 
11 1 4 5 6 41 42 43 34 35 27 28 
11 1 4 5 6 41 42 43 34 35 20 21 
12 1 4 5 6 41 41 42 43 7 8 9 10 
10 1 4 5 6 41 41 42 43 27 28 
11 1 4 5 6 41 41 41 7 8 9 10 
11 1 4 5 6 41 41 41 7 15 9 17 
9 1 4 5 6 41 41 41 27 28 
12 1 4 5 6 41 41 44 45 7 8 9 10 
10 1 4 5 6 41 41 44 45 27 28 
12 1 4 5 6 36 37 11 12 13 14 27 28 
12 1 4 5 6 41 41 30 31 7 8 9 10 
12 1 4 5 6 41 41 30 31 7 15 9 17 
10 1 4 5 6 41 41 30 31 27 28 
13 1 4 5 6 41 41 30 31 29 7 20 9 21 
12 1 4 5 6 41 41 46 47 7 8 9 10 
10 1 4 5 6 41 41 46 47 27 28 
13 1 4 5 6 41 41 46 47 29 7 20 9 21 
12 1 4 5 6 41 41 27 28 7 8 9 10 
12 1 4 5 6 41 41 27 28 7 15 9 17 
10 1 4 5 6 41 41 27 28 27 28 
8 1 4 5 6 7 8 9 10 
12 1 4 5 6 36 37 11 12 13 14 20 21 
11 1 4 5 6 41 41 33 7 8 9 10 
9 1 4 5 6 41 41 33 27 28 
12 1 4 5 6 41 41 38 39 7 8 9 10 
12 1 4 5 6 41 41 38 39 7 15 9 17 
10 1 4 5 6 41 41 38 39 27 28 
11 1 4 5 6 41 41 40 7 8 9 10 
9 1 4 5 6 41 41 40 27 28 
13 1 4 5 6 41 44 45 42 43 7 8 9 10 
11 1 4 5 6 41 44 45 42 43 27 28 
15 1 4 5 6 41 44 45 11 12 13 14 7 8 9 10 
10 1 4 5 6 36 37 7 8 9 10 
14 1 4 5 6 41 44 45 11 12 13 14 15 16 17 
13 1 4 5 6 41 44 45 11 12 13 14 27 28 
13 1 4 5 6 41 44 45 11 12 13 14 20 21 
13 1 4 5 6 41 44 45 44 45 7 8 9 10 
11 1 4 5 6 41 44 45 44 45 27 28 
16 1 4 5 6 41 44 45 22 29 7 23 25 7 8 9 10 
16 1 4 5 6 41 44 45 22 29 7 23 25 7 15 9 17 
14 1 4 5 6 41 44 45 22 29 7 23 25 27 28 
13 1 4 5 6 41 44 45 27 28 7 8 9 10 
13 1 4 5 6 41 44 45 27 28 7 15 9 17 
10 1 4 5 6 36 37 7 8 9 10 
11 1 4 5 6 41 44 45 27 28 27 28 
13 1 4 5 6 41 44 45 34 35 7 8 9 10 
12 1 4 5 6 41 44 45 34 35 15 16 17 
11 1 4 5 6 41 44 45 34 35 27 28 
11 1 4 5 6 41 44 45 34 35 20 21 
13 1 4 5 6 41 30 31 42 43 7 8 9 10 
11 1 4 5 6 41 30 31 42 43 27 28 
13 1 4 5 6 41 30 31 44 45 7 8 9 10 
11 1 4 5 6 41 30 31 44 45 27 28 
13 1 4 5 6 41 30 31 30 31 7 8 9 10 
10 1 4 5 6 36 37 7 8 9 10 
13 1 4 5 6 41 30 31 30 31 7 15 9 17 
11 1 4 5 6 41 30 31 30 31 27 28 
14 1 4 5 6 41 30 31 30 31 29 7 20 9 21 
13 1 4 5 6 41 30 31 46 47 7 8 9 10 
11 1 4 5 6 41 30 31 46 47 27 28 
14 1 4 5 6 41 30 31 46 47 29 7 20 9 21 
16 1 4 5 6 41 30 31 22 29 7 23 25 7 8 9 10 
16 1 4 5 6 41 30 31 22 29 7 23 25 7 15 9 17 
14 1 4 5 6 41 30 31 22 29 7 23 25 27 28 
13 1 4 5 6 41 30 31 27 28 7 8 9 10 
10 1 4 5 6 36 37 7 8 9 10 
13 1 4 5 6 41 30 31 27 28 7 15 9 17 
11 1 4 5 6 41 30 31 27 28 27 28 
12 1 4 5 6 41 30 31 33 7 8 9 10 
10 1 4 5 6 41 30 31 33 27 28 
12 1 4 5 6 41 30 31 40 7 8 9 10 
10 1 4 5 6 41 30 31 40 27 28 
13 1 4 5 6 41 46 47 42 43 7 8 9 10 
11 1 4 5 6 41 46 47 42 43 27 28 
15 1 4 5 6 41 46 47 11 12 13 14 7 8 9 10 
14 1 4 5 6 41 46 47 11 12 13 14 15 16 17 
11 1 4 5 6 36 37 41 7 8 9 10 
13 1 4 5 6 41 46 47 11 12 13 14 27 28 
13 1 4 5 6 41 46 47 11 12 13 14 20 21 
13 1 4 5 6 41 46 47 44 45 7 8 9 10 
11 1 4 5 6 41 46 47 44 45 27 28 
13 1 4 5 6 41 46 47 46 47 7 8 9 10 
11 1 4 5 6 41 46 47 46 47 27 28 
14 1 4 5 6 41 46 47 46 47 29 7 20 9 21 
16 1 4 5 6 41 46 47 22 29 7 23 25 7 8 9 10 
16 1 4 5 6 41 46 47 22 29 7 23 25 7 15 9 17 
14 1 4 5 6 41 46 47 22 29 7 23 25 27 28 
10 1 4 5 6 36 37 41 15 16 17 
13 1 4 5 6 41 46 47 27 28 7 8 9 10 
13 1 4 5 6 41 46 47 27 28 7 15 9 17 
11 1 4 5 6 41 46 47 27 28 27 28 
13 1 4 5 6 41 46 47 34 35 7 8 9 10 
12 1 4 5 6 41 46 47 34 35 15 16 17 
11 1 4 5 6 41 46 47 34 35 27 28 
11 1 4 5 6 41 46 47 34 35 20 21 
12 1 4 5 6 41 46 47 40 7 8 9 10 
10 1 4 5 6 41 46 47 40 27 28 
13 1 4 5 6 41 27 28 30 31 7 8 9 10 
9 1 4 5 6 36 37 41 27 28 
13 1 4 5 6 41 27 28 30 31 7 15 9 17 
11 1 4 5 6 41 27 28 30 31 27 28 
14 1 4 5 6 41 27 28 30 31 29 7 20 9 21 
13 1 4 5 6 41 27 28 27 28 7 8 9 10 
13 1 4 5 6 41 27 28 27 28 7 15 9 17 
11 1 4 5 6 41 27 28 27 28 27 28 
13 1 4 5 6 41 27 28 38 39 7 8 9 10 
13 1 4 5 6 41 27 28 38 39 7 15 9 17 
11 1 4 5 6 41 27 28 38 39 27 28 
12 1 4 5 6 41 33 42 43 7 8 9 10 
12 1 4 5 6 36 37 41 29 7 20 9 21 
10 1 4 5 6 41 33 42 43 27 28 
12 1 4 5 6 41 33 44 45 7 8 9 10 
10 1 4 5 6 41 33 44 45 27 28 
12 1 4 5 6 41 33 46 47 7 8 9 10 
10 1 4 5 6 41 33 46 47 27 28 
13 1 4 5 6 41 33 46 47 29 7 20 9 21 
12 1 4 5 6 41 33 27 28 7 8 9 10 
12 1 4 5 6 41 33 27 28 7 15 9 17 
10 1 4 5 6 41 33 27 28 27 28 
11 1 4 5 6 41 33 33 7 8 9 10 
12 1 4 5 6 36 37 44 45 7 8 9 10 
9 1 4 5 6 41 33 33 27 28 
11 1 4 5 6 41 33 40 7 8 9 10 
9 1 4 5 6 41 33 40 27 28 
13 1 4 5 6 41 38 39 42 43 7 8 9 10 
11 1 4 5 6 41 38 39 42 43 27 28 
13 1 4 5 6 41 38 39 44 45 7 8 9 10 
11 1 4 5 6 41 38 39 44 45 27 28 
13 1 4 5 6 41 38 39 30 31 7 8 9 10 
13 1 4 5 6 41 38 39 30 31 7 15 9 17 
11 1 4 5 6 41 38 39 30 31 27 28 
9 1 4 5 6 41 7 8 9 10 
11 1 4 5 6 36 37 44 45 15 16 17 
14 1 4 5 6 41 38 39 30 31 29 7 20 9 21 
13 1 4 5 6 41 38 39 46 47 7 8 9 10 
11 1 4 5 6 41 38 39 46 47 27 28 
14 1 4 5 6 41 38 39 46 47 29 7 20 9 21 
16 1 4 5 6 41 38 39 22 29 7 23 25 7 8 9 10 
16 1 4 5 6 41 38 39 22 29 7 23 25 7 15 9 17 
14 1 4 5 6 41 38 39 22 29 7 23 25 27 28 
13 1 4 5 6 41 38 39 27 28 7 8 9 10 
13 1 4 5 6 41 38 39 27 28 7 15 9 17 
11 1 4 5 6 41 38 39 27 28 27 28 
10 1 4 5 6 36 37 44 45 27 28 
12 1 4 5 6 41 38 39 33 7 8 9 10 
10 1 4 5 6 41 38 39 33 27 28 
13 1 4 5 6 41 38 39 38 39 7 8 9 10 
13 1 4 5 6 41 38 39 38 39 7 15 9 17 
11 1 4 5 6 41 38 39 38 39 27 28 
12 1 4 5 6 41 38 39 40 7 8 9 10 
10 1 4 5 6 41 38 39 40 27 28 
12 1 4 5 6 41 40 42 43 7 8 9 10 
10 1 4 5 6 41 40 42 43 27 28 
12 1 4 5 6 41 40 44 45 7 8 9 10 
13 1 4 5 6 36 37 44 45 29 7 20 9 21 
10 1 4 5 6 41 40 44 45 27 28 
12 1 4 5 6 41 40 27 28 7 8 9 10 
12 1 4 5 6 41 40 27 28 7 15 9 17 
10 1 4 5 6 41 40 27 28 27 28 
11 1 4 5 6 41 40 40 7 8 9 10 
9 1 4 5 6 41 40 40 27 28 
14 1 4 5 6 44 45 42 43 42 43 7 8 9 10 
12 1 4 5 6 44 45 42 43 42 43 27 28 
16 1 4 5 6 44 45 42 43 11 12 13 14 7 8 9 10 
15 1 4 5 6 44 45 42 43 11 12 13 14 15 16 17 
12 1 4 5 6 36 37 18 19 7 8 9 10 
14 1 4 5 6 44 45 42 43 11 12 13 14 27 28 
14 1 4 5 6 44 45 42 43 11 12 13 14 20 21 
17 1 4 5 6 44 45 42 43 22 29 7 23 25 7 8 9 10 
17 1 4 5 6 44 45 42 43 22 29 7 23 25 7 15 9 17 
15 1 4 5 6 44 45 42 43 22 29 7 23 25 27 28 
14 1 4 5 6 44 45 42 43 27 28 7 8 9 10 
14 1 4 5 6 44 45 42 43 27 28 7 15 9 17 
12 1 4 5 6 44 45 42 43 27 28 27 28 
14 1 4 5 6 44 45 42 43 34 35 7 8 9 10 
13 1 4 5 6 44 45 42 43 34 35 15 16 17 
11 1 4 5 6 36 37 18 19 15 16 17 
12 1 4 5 6 44 45 42 43 34 35 27 28 
12 1 4 5 6 44 45 42 43 34 35 20 21 
16 1 4 5 6 44 45 11 12 13 14 42 43 7 8 9 10 
14 1 4 5 6 44 45 11 12 13 14 42 43 27 28 
18 1 4 5 6 44 45 11 12 13 14 11 12 13 14 7 8 9 10 
17 1 4 5 6 44 45 11 12 13 14 11 12 13 14 15 16 17 
16 1 4 5 6 44 45 11 12 13 14 11 12 13 14 27 28 
16 1 4 5 6 44 45 11 12 13 14 11 12 13 14 20 21 
15 1 4 5 6 44 45 11 12 13 14 41 7 8 9 10 
14 1 4 5 6 44 45 11 12 13 14 41 15 16 17 
10 1 4 5 6 36 37 18 19 27 28 
13 1 4 5 6 44 45 11 12 13 14 41 27 28 
16 1 4 5 6 44 45 11 12 13 14 44 45 7 8 9 10 
14 1 4 5 6 44 45 11 12 13 14 44 45 27 28 
16 1 4 5 6 44 45 11 12 13 14 18 19 7 8 9 10 
15 1 4 5 6 44 45 11 12 13 14 18 19 15 16 17 
14 1 4 5 6 44 45 11 12 13 14 18 19 27 28 
14 1 4 5 6 44 45 11 12 13 14 18 19 20 21 
16 1 4 5 6 44 45 11 12 13 14 30 31 7 8 9 10 
15 1 4 5 6 44 45 11 12 13 14 30 31 15 16 17 
14 1 4 5 6 44 45 11 12 13 14 30 31 27 28 
13 1 4 5 6 36 37 18 19 29 7 20 9 21 
14 1 4 5 6 44 45 11 12 13 14 30 31 20 21 
16 1 4 5 6 44 45 11 12 13 14 46 47 7 8 9 10 
14 1 4 5 6 44 45 11 12 13 14 46 47 27 28 
14 1 4 5 6 44 45 11 12 13 14 46 47 20 21 
19 1 4 5 6 44 45 11 12 13 14 22 23 26 24 25 7 8 9 10 
18 1 4 5 6 44 45 11 12 13 14 22 23 24 25 7 8 9 10 
18 1 4 5 6 44 45 11 12 13 14 22 23 26 24 25 15 16 17 
17 1 4 5 6 44 45 11 12 13 14 22 23 24 25 15 16 17 
17 1 4 5 6 44 45 11 12 13 14 22 23 26 24 25 27 28 
16 1 4 5 6 44 45 11 12 13 14 22 23 24 25 27 28 
12 1 4 5 6 36 37 30 31 7 8 9 10 
15 1 4 5 6 44 45 11 12 13 14 15 16 17 8 10 
16 1 4 5 6 44 45 11 12 13 14 15 16 17 15 16 17 
17 1 4 5 6 44 45 11 12 13 14 15 16 17 7 27 9 28 
18 1 4 5 6 44 45 11 12 13 14 15 16 17 29 7 20 9 21 
16 1 4 5 6 44 45 11 12 13 14 27 28 7 8 9 10 
15 1 4 5 6 44 45 11 12 13 14 27 28 15 16 17 
14 1 4 5 6 44 45 11 12 13 14 27 28 27 28 
16 1 4 5 6 44 45 11 12 13 14 13 32 7 8 9 10 
15 1 4 5 6 44 45 11 12 13 14 13 32 15 16 17 
14 1 4 5 6 44 45 11 12 13 14 13 32 27 28 
11 1 4 5 6 36 37 30 31 15 16 17 
15 1 4 5 6 44 45 11 12 13 14 33 7 8 9 10 
13 1 4 5 6 44 45 11 12 13 14 33 27 28 
16 1 4 5 6 44 45 11 12 13 14 34 35 7 8 9 10 
15 1 4 5 6 44 45 11 12 13 14 34 35 15 16 17 
14 1 4 5 6 44 45 11 12 13 14 34 35 27 28 
14 1 4 5 6 44 45 11 12 13 14 34 35 20 21 
16 1 4 5 6 44 45 11 12 13 14 36 37 7 8 9 10 
15 1 4 5 6 44 45 11 12 13 14 36 37 15 16 17 
14 1 4 5 6 44 45 11 12 13 14 36 37 27 28 
14 1 4 5 6 44 45 11 12 13 14 36 37 20 21 
10 1 4 5 6 36 37 30 31 27 28 
16 1 4 5 6 44 45 11 12 13 14 38 39 7 8 9 10 
15 1 4 5 6 44 45 11 12 13 14 38 39 15 16 17 
14 1 4 5 6 44 45 11 12 13 14 38 39 27 28 
15 1 4 5 6 44 45 11 12 13 14 40 7 8 9 10 
13 1 4 5 6 44 45 11 12 13 14 40 27 28 
16 1 4 5 6 44 45 11 12 13 14 20 21 7 8 9 10 
15 1 4 5 6 44 45 11 12 13 14 20 21 15 16 17 
14 1 4 5 6 44 45 11 12 13 14 20 21 27 28 
14 1 4 5 6 44 45 11 12 13 14 20 21 20 21 
14 1 4 5 6 44 45 44 45 42 43 7 8 9 10 
9 1 4 5 6 41 7 15 9 17 
13 1 4 5 6 36 37 30 31 29 7 20 9 21 
12 1 4 5 6 44 45 44 45 42 43 27 28 
16 1 4 5 6 44 45 44 45 11 12 13 14 7 8 9 10 
15 1 4 5 6 44 45 44 45 11 12 13 14 15 16 17 
14 1 4 5 6 44 45 44 45 11 12 13 14 27 28 
14 1 4 5 6 44 45 44 45 11 12 13 14 20 21 
14 1 4 5 6 44 45 44 45 44 45 7 8 9 10 
12 1 4 5 6 44 45 44 45 44 45 27 28 
17 1 4 5 6 44 45 44 45 22 29 7 23 25 7 8 9 10 
17 1 4 5 6 44 45 44 45 22 29 7 23 25 7 15 9 17 
15 1 4 5 6 44 45 44 45 22 29 7 23 25 27 28 
12 1 4 5 6 36 37 46 47 7 8 9 10 
14 1 4 5 6 44 45 44 45 27 28 7 8 9 10 
14 1 4 5 6 44 45 44 45 27 28 7 15 9 17 
12 1 4 5 6 44 45 44 45 27 28 27 28 
14 1 4 5 6 44 45 44 45 34 35 7 8 9 10 
13 1 4 5 6 44 45 44 45 34 35 15 16 17 
12 1 4 5 6 44 45 44 45 34 35 27 28 
12 1 4 5 6 44 45 44 45 34 35 20 21 
17 1 4 5 6 44 45 22 29 7 23 25 42 43 7 8 9 10 
15 1 4 5 6 44 45 22 29 7 23 25 42 43 27 28 
19 1 4 5 6 44 45 22 29 7 23 25 11 12 13 14 7 8 9 10 
11 1 4 5 6 36 37 46 47 15 16 17 
18 1 4 5 6 44 45 22 29 7 23 25 11 12 13 14 15 16 17 
17 1 4 5 6 44 45 22 29 7 23 25 11 12 13 14 27 28 
17 1 4 5 6 44 45 22 29 7 23 25 11 12 13 14 20 21 
16 1 4 5 6 44 45 22 29 7 23 25 41 7 8 9 10 
16 1 4 5 6 44 45 22 29 7 23 25 41 7 15 9 17 
14 1 4 5 6 44 45 22 29 7 23 25 41 27 28 
17 1 4 5 6 44 45 22 29 7 23 25 44 45 7 8 9 10 
15 1 4 5 6 44 45 22 29 7 23 25 44 45 27 28 
17 1 4 5 6 44 45 22 29 7 23 25 18 19 7 8 9 10 
17 1 4 5 6 44 45 22 29 7 23 25 18 19 7 15 9 17 
10 1 4 5 6 36 37 46 47 27 28 
15 1 4 5 6 44 45 22 29 7 23 25 18 19 27 28 
18 1 4 5 6 44 45 22 29 7 23 25 18 19 29 7 20 9 21 
17 1 4 5 6 44 45 22 29 7 23 25 30 31 7 8 9 10 
17 1 4 5 6 44 45 22 29 7 23 25 30 31 7 15 9 17 
15 1 4 5 6 44 45 22 29 7 23 25 30 31 27 28 
18 1 4 5 6 44 45 22 29 7 23 25 30 31 29 7 20 9 21 
17 1 4 5 6 44 45 22 29 7 23 25 46 47 7 8 9 10 
15 1 4 5 6 44 45 22 29 7 23 25 46 47 27 28 
18 1 4 5 6 44 45 22 29 7 23 25 46 47 29 7 20 9 21 
20 1 4 5 6 44 45 22 29 7 23 25 22 29 7 23 25 7 8 9 10 
10 1 4 5 6 36 37 46 47 20 21 
20 1 4 5 6 44 45 22 29 7 23 25 22 29 7 23 25 7 15 9 17 
18 1 4 5 6 44 45 22 29 7 23 25 22 29 7 23 25 27 28 
17 1 4 5 6 44 45 22 29 7 23 25 27 28 7 8 9 10 
17 1 4 5 6 44 45 22 29 7 23 25 27 28 7 15 9 17 
15 1 4 5 6 44 45 22 29 7 23 25 27 28 27 28 
17 1 4 5 6 44 45 22 29 7 23 25 13 32 7 8 9 10 
17 1 4 5 6 44 45 22 29 7 23 25 13 32 7 15 9 17 
15 1 4 5 6 44 45 22 29 7 23 25 13 32 27 28 
16 1 4 5 6 44 45 22 29 7 23 25 33 7 8 9 10 
14 1 4 5 6 44 45 22 29 7 23 25 33 27 28 
15 1 4 5 6 36 37 22 29 7 23 25 7 8 9 10 
17 1 4 5 6 44 45 22 29 7 23 25 34 35 7 8 9 10 
16 1 4 5 6 44 45 22 29 7 23 25 34 35 15 16 17 
15 1 4 5 6 44 45 22 29 7 23 25 34 35 27 28 
15 1 4 5 6 44 45 22 29 7 23 25 34 35 20 21 
17 1 4 5 6 44 45 22 29 7 23 25 36 37 7 8 9 10 
16 1 4 5 6 44 45 22 29 7 23 25 36 37 15 16 17 
15 1 4 5 6 44 45 22 29 7 23 25 36 37 27 28 
18 1 4 5 6 44 45 22 29 7 23 25 36 37 29 7 20 9 21 
17 1 4 5 6 44 45 22 29 7 23 25 38 39 7 8 9 10 
17 1 4 5 6 44 45 22 29 7 23 25 38 39 7 15 9 17 
14 1 4 5 6 36 37 22 29 7 23 25 15 16 17 
15 1 4 5 6 44 45 22 29 7 23 25 38 39 27 28 
16 1 4 5 6 44 45 22 29 7 23 25 40 7 8 9 10 
14 1 4 5 6 44 45 22 29 7 23 25 40 27 28 
14 1 4 5 6 44 45 27 28 30 31 7 8 9 10 
14 1 4 5 6 44 45 27 28 30 31 7 15 9 17 
12 1 4 5 6 44 45 27 28 30 31 27 28 
15 1 4 5 6 44 45 27 28 30 31 29 7 20 9 21 
14 1 4 5 6 44 45 27 28 27 28 7 8 9 10 
14 1 4 5 6 44 45 27 28 27 28 7 15 9 17 
12 1 4 5 6 44 45 27 28 27 28 27 28 
13 1 4 5 6 36 37 22 29 7 23 25 27 28 
14 1 4 5 6 44 45 27 28 38 39 7 8 9 10 
14 1 4 5 6 44 45 27 28 38 39 7 15 9 17 
12 1 4 5 6 44 45 27 28 38 39 27 28 
14 1 4 5 6 44 45 34 35 42 43 7 8 9 10 
12 1 4 5 6 44 45 34 35 42 43 27 28 
16 1 4 5 6 44 45 34 35 11 12 13 14 7 8 9 10 
15 1 4 5 6 44 45 34 35 11 12 13 14 15 16 17 
14 1 4 5 6 44 45 34 35 11 12 13 14 27 28 
14 1 4 5 6 44 45 34 35 11 12 13 14 20 21 
13 1 4 5 6 44 45 34 35 41 7 8 9 10 
16 1 4 5 6 36 37 22 29 7 23 25 29 7 20 9 21 
12 1 4 5 6 44 45 34 35 41 15 16 17 
11 1 4 5 6 44 45 34 35 41 27 28 
14 1 4 5 6 44 45 34 35 44 45 7 8 9 10 
12 1 4 5 6 44 45 34 35 44 45 27 28 
14 1 4 5 6 44 45 34 35 18 19 7 8 9 10 
13 1 4 5 6 44 45 34 35 18 19 15 16 17 
12 1 4 5 6 44 45 34 35 18 19 27 28 
12 1 4 5 6 44 45 34 35 18 19 20 21 
14 1 4 5 6 44 45 34 35 30 31 7 8 9 10 
13 1 4 5 6 44 45 34 35 30 31 15 16 17 
11 1 4 5 6 36 37 15 16 17 8 10 
12 1 4 5 6 44 45 34 35 30 31 27 28 
12 1 4 5 6 44 45 34 35 30 31 20 21 
14 1 4 5 6 44 45 34 35 46 47 7 8 9 10 
12 1 4 5 6 44 45 34 35 46 47 27 28 
12 1 4 5 6 44 45 34 35 46 47 20 21 
17 1 4 5 6 44 45 34 35 22 23 26 24 25 7 8 9 10 
16 1 4 5 6 44 45 34 35 22 23 24 25 7 8 9 10 
16 1 4 5 6 44 45 34 35 22 23 26 24 25 15 16 17 
15 1 4 5 6 44 45 34 35 22 23 24 25 15 16 17 
15 1 4 5 6 44 45 34 35 22 23 26 24 25 27 28 
7 1 4 5 6 41 27 28 
12 1 4 5 6 36 37 15 16 17 15 16 17 
14 1 4 5 6 44 45 34 35 22 23 24 25 27 28 
13 1 4 5 6 44 45 34 35 15 16 17 8 10 
14 1 4 5 6 44 45 34 35 15 16 17 15 16 17 
15 1 4 5 6 44 45 34 35 15 16 17 7 27 9 28 
16 1 4 5 6 44 45 34 35 15 16 17 29 7 20 9 21 
14 1 4 5 6 44 45 34 35 27 28 7 8 9 10 
13 1 4 5 6 44 45 34 35 27 28 15 16 17 
12 1 4 5 6 44 45 34 35 27 28 27 28 
14 1 4 5 6 44 45 34 35 13 32 7 8 9 10 
13 1 4 5 6 44 45 34 35 13 32 15 16 17 
13 1 4 5 6 36 37 15 16 17 7 27 9 28 
12 1 4 5 6 44 45 34 35 13 32 27 28 
13 1 4 5 6 44 45 34 35 33 7 8 9 10 
11 1 4 5 6 44 45 34 35 33 27 28 
14 1 4 5 6 44 45 34 35 34 35 7 8 9 10 
13 1 4 5 6 44 45 34 35 34 35 15 16 17 
12 1 4 5 6 44 45 34 35 34 35 27 28 
12 1 4 5 6 44 45 34 35 34 35 20 21 
14 1 4 5 6 44 45 34 35 36 37 7 8 9 10 
13 1 4 5 6 44 45 34 35 36 37 15 16 17 
12 1 4 5 6 44 45 34 35 36 37 27 28 
14 1 4 5 6 36 37 15 16 17 29 7 20 9 21 
12 1 4 5 6 44 45 34 35 36 37 20 21 
14 1 4 5 6 44 45 34 35 38 39 7 8 9 10 
13 1 4 5 6 44 45 34 35 38 39 15 16 17 
12 1 4 5 6 44 45 34 35 38 39 27 28 
13 1 4 5 6 44 45 34 35 40 7 8 9 10 
11 1 4 5 6 44 45 34 35 40 27 28 
14 1 4 5 6 44 45 34 35 20 21 7 8 9 10 
13 1 4 5 6 44 45 34 35 20 21 15 16 17 
12 1 4 5 6 44 45 34 35 20 21 27 28 
12 1 4 5 6 44 45 34 35 20 21 20 21 
12 1 4 5 6 36 37 27 28 7 8 9 10 
14 1 4 5 6 18 19 42 43 42 43 7 8 9 10 
12 1 4 5 6 18 19 42 43 42 43 27 28 
16 1 4 5 6 18 19 42 43 11 12 13 14 7 8 9 10 
15 1 4 5 6 18 19 42 43 11 12 13 14 15 16 17 
14 1 4 5 6 18 19 42 43 11 12 13 14 27 28 
14 1 4 5 6 18 19 42 43 11 12 13 14 20 21 
17 1 4 5 6 18 19 42 43 22 29 7 23 25 7 8 9 10 
17 1 4 5 6 18 19 42 43 22 29 7 23 25 7 15 9 17 
15 1 4 5 6 18 19 42 43 22 29 7 23 25 27 28 
14 1 4 5 6 18 19 42 43 27 28 7 8 9 10 
11 1 4 5 6 36 37 27 28 15 16 17 
14 1 4 5 6 18 19 42 43 27 28 7 15 9 17 
12 1 4 5 6 18 19 42 43 27 28 27 28 
14 1 4 5 6 18 19 42 43 34 35 7 8 9 10 
13 1 4 5 6 18 19 42 43 34 35 15 16 17 
12 1 4 5 6 18 19 42 43 34 35 27 28 
12 1 4 5 6 18 19 42 43 34 35 20 21 
13 1 4 5 6 18 19 41 42 43 7 8 9 10 
11 1 4 5 6 18 19 41 42 43 27 28 
12 1 4 5 6 18 19 41 41 7 8 9 10 
12 1 4 5 6 18 19 41 41 7 15 9 17 
10 1 4 5 6 36 37 27 28 27 28 
10 1 4 5 6 18 19 41 41 27 28 
13 1 4 5 6 18 19 41 44 45 7 8 9 10 
11 1 4 5 6 18 19 41 44 45 27 28 
13 1 4 5 6 18 19 41 30 31 7 8 9 10 
13 1 4 5 6 18 19 41 30 31 7 15 9 17 
11 1 4 5 6 18 19 41 30 31 27 28 
14 1 4 5 6 18 19 41 30 31 29 7 20 9 21 
13 1 4 5 6 18 19 41 46 47 7 8 9 10 
11 1 4 5 6 18 19 41 46 47 27 28 
14 1 4 5 6 18 19 41 46 47 29 7 20 9 21 
13 1 4 5 6 36 37 27 28 29 7 20 9 21 
13 1 4 5 6 18 19 41 27 28 7 8 9 10 
13 1 4 5 6 18 19 41 27 28 7 15 9 17 
11 1 4 5 6 18 19 41 27 28 27 28 
12 1 4 5 6 18 19 41 33 7 8 9 10 
10 1 4 5 6 18 19 41 33 27 28 
13 1 4 5 6 18 19 41 38 39 7 8 9 10 
13 1 4 5 6 18 19 41 38 39 7 15 9 17 
11 1 4 5 6 18 19 41 38 39 27 28 
12 1 4 5 6 18 19 41 40 7 8 9 10 
10 1 4 5 6 18 19 41 40 27 28 
12 1 4 5 6 36 37 13 32 7 8 9 10 
14 1 4 5 6 18 19 44 45 42 43 7 8 9 10 
12 1 4 5 6 18 19 44 45 42 43 27 28 
16 1 4 5 6 18 19 44 45 11 12 13 14 7 8 9 10 
15 1 4 5 6 18 19 44 45 11 12 13 14 15 16 17 
14 1 4 5 6 18 19 44 45 11 12 13 14 27 28 
14 1 4 5 6 18 19 44 45 11 12 13 14 20 21 
14 1 4 5 6 18 19 44 45 44 45 7 8 9 10 
12 1 4 5 6 18 19 44 45 44 45 27 28 
17 1 4 5 6 18 19 44 45 22 29 7 23 25 7 8 9 10 
17 1 4 5 6 18 19 44 45 22 29 7 23 25 7 15 9 17 
11 1 4 5 6 36 37 13 32 15 16 17 
15 1 4 5 6 18 19 44 45 22 29 7 23 25 27 28 
14 1 4 5 6 18 19 44 45 27 28 7 8 9 10 
14 1 4 5 6 18 19 44 45 27 28 7 15 9 17 
12 1 4 5 6 18 19 44 45 27 28 27 28 
14 1 4 5 6 18 19 44 45 34 35 7 8 9 10 
13 1 4 5 6 18 19 44 45 34 35 15 16 17 
12 1 4 5 6 18 19 44 45 34 35 27 28 
12 1 4 5 6 18 19 44 45 34 35 20 21 
14 1 4 5 6 18 19 18 19 42 43 7 8 9 10 
12 1 4 5 6 18 19 18 19 42 43 27 28 
10 1 4 5 6 36 37 13 32 27 28 
13 1 4 5 6 18 19 18 19 41 7 8 9 10 
13 1 4 5 6 18 19 18 19 41 7 15 9 17 
11 1 4 5 6 18 19 18 19 41 27 28 
14 1 4 5 6 18 19 18 19 44 45 7 8 9 10 
12 1 4 5 6 18 19 18 19 44 45 27 28 
14 1 4 5 6 18 19 18 19 18 19 7 8 9 10 
14 1 4 5 6 18 19 18 19 18 19 7 15 9 17 
12 1 4 5 6 18 19 18 19 18 19 27 28 
15 1 4 5 6 18 19 18 19 18 19 29 7 20 9 21 
14 1 4 5 6 18 19 18 19 30 31 7 8 9 10 
8 1 4 5 6 7 15 9 17 
10 1 4 5 6 41 29 7 20 9 21 
13 1 4 5 6 36 37 13 32 29 7 20 9 21 
14 1 4 5 6 18 19 18 19 30 31 7 15 9 17 
12 1 4 5 6 18 19 18 19 30 31 27 28 
15 1 4 5 6 18 19 18 19 30 31 29 7 20 9 21 
14 1 4 5 6 18 19 18 19 46 47 7 8 9 10 
12 1 4 5 6 18 19 18 19 46 47 27 28 
15 1 4 5 6 18 19 18 19 46 47 29 7 20 9 21 
17 1 4 5 6 18 19 18 19 22 29 7 23 25 7 8 9 10 
17 1 4 5 6 18 19 18 19 22 29 7 23 25 7 15 9 17 
15 1 4 5 6 18 19 18 19 22 29 7 23 25 27 28 
14 1 4 5 6 18 19 18 19 27 28 7 8 9 10 
11 1 4 5 6 36 37 33 7 8 9 10 
14 1 4 5 6 18 19 18 19 27 28 7 15 9 17 
12 1 4 5 6 18 19 18 19 27 28 27 28 
14 1 4 5 6 18 19 18 19 13 32 7 8 9 10 
14 1 4 5 6 18 19 18 19 13 32 7 15 9 17 
12 1 4 5 6 18 19 18 19 13 32 27 28 
13 1 4 5 6 18 19 18 19 33 7 8 9 10 
11 1 4 5 6 18 19 18 19 33 27 28 
14 1 4 5 6 18 19 18 19 36 37 7 8 9 10 
13 1 4 5 6 18 19 18 19 36 37 15 16 17 
12 1 4 5 6 18 19 18 19 36 37 27 28 
10 1 4 5 6 36 37 33 15 16 17 
15 1 4 5 6 18 19 18 19 36 37 29 7 20 9 21 
14 1 4 5 6 18 19 18 19 38 39 7 8 9 10 
14 1 4 5 6 18 19 18 19 38 39 7 15 9 17 
12 1 4 5 6 18 19 18 19 38 39 27 28 
13 1 4 5 6 18 19 18 19 40 7 8 9 10 
11 1 4 5 6 18 19 18 19 40 27 28 
14 1 4 5 6 18 19 30 31 42 43 7 8 9 10 
12 1 4 5 6 18 19 30 31 42 43 27 28 
14 1 4 5 6 18 19 30 31 44 45 7 8 9 10 
12 1 4 5 6 18 19 30 31 44 45 27 28 
9 1 4 5 6 36 37 33 27 28 
14 1 4 5 6 18 19 30 31 30 31 7 8 9 10 
14 1 4 5 6 18 19 30 31 30 31 7 15 9 17 
12 1 4 5 6 18 19 30 31 30 31 27 28 
15 1 4 5 6 18 19 30 31 30 31 29 7 20 9 21 
14 1 4 5 6 18 19 30 31 46 47 7 8 9 10 
12 1 4 5 6 18 19 30 31 46 47 27 28 
15 1 4 5 6 18 19 30 31 46 47 29 7 20 9 21 
17 1 4 5 6 18 19 30 31 22 29 7 23 25 7 8 9 10 
17 1 4 5 6 18 19 30 31 22 29 7 23 25 7 15 9 17 
15 1 4 5 6 18 19 30 31 22 29 7 23 25 27 28 
12 1 4 5 6 36 37 33 29 7 20 9 21 
14 1 4 5 6 18 19 30 31 27 28 7 8 9 10 
14 1 4 5 6 18 19 30 31 27 28 7 15 9 17 
12 1 4 5 6 18 19 30 31 27 28 27 28 
13 1 4 5 6 18 19 30 31 33 7 8 9 10 
11 1 4 5 6 18 19 30 31 33 27 28 
13 1 4 5 6 18 19 30 31 40 7 8 9 10 
11 1 4 5 6 18 19 30 31 40 27 28 
14 1 4 5 6 18 19 46 47 42 43 7 8 9 10 
12 1 4 5 6 18 19 46 47 42 43 27 28 
16 1 4 5 6 18 19 46 47 11 12 13 14 7 8 9 10 
12 1 4 5 6 36 37 34 35 7 8 9 10 
15 1 4 5 6 18 19 46 47 11 12 13 14 15 16 17 
14 1 4 5 6 18 19 46 47 11 12 13 14 27 28 
14 1 4 5 6 18 19 46 47 11 12 13 14 20 21 
14 1 4 5 6 18 19 46 47 44 45 7 8 9 10 
12 1 4 5 6 18 19 46 47 44 45 27 28 
14 1 4 5 6 18 19 46 47 46 47 7 8 9 10 
12 1 4 5 6 18 19 46 47 46 47 27 28 
15 1 4 5 6 18 19 46 47 46 47 29 7 20 9 21 
17 1 4 5 6 18 19 46 47 22 29 7 23 25 7 8 9 10 
17 1 4 5 6 18 19 46 47 22 29 7 23 25 7 15 9 17 
11 1 4 5 6 36 37 34 35 15 16 17 
15 1 4 5 6 18 19 46 47 22 29 7 23 25 27 28 
14 1 4 5 6 18 19 46 47 27 28 7 8 9 10 
14 1 4 5 6 18 19 46 47 27 28 7 15 9 17 
12 1 4 5 6 18 19 46 47 27 28 27 28 
14 1 4 5 6 18 19 46 47 34 35 7 8 9 10 
13 1 4 5 6 18 19 46 47 34 35 15 16 17 
12 1 4 5 6 18 19 46 47 34 35 27 28 
12 1 4 5 6 18 19 46 47 34 35 20 21 
13 1 4 5 6 18 19 46 47 40 7 8 9 10 
11 1 4 5 6 18 19 46 47 40 27 28 
10 1 4 5 6 36 37 34 35 27 28 
17 1 4 5 6 18 19 22 29 7 23 25 42 43 7 8 9 10 
15 1 4 5 6 18 19 22 29 7 23 25 42 43 27 28 
19 1 4 5 6 18 19 22 29 7 23 25 11 12 13 14 7 8 9 10 
18 1 4 5 6 18 19 22 29 7 23 25 11 12 13 14 15 16 17 
17 1 4 5 6 18 19 22 29 7 23 25 11 12 13 14 27 28 
17 1 4 5 6 18 19 22 29 7 23 25 11 12 13 14 20 21 
16 1 4 5 6 18 19 22 29 7 23 25 41 7 8 9 10 
16 1 4 5 6 18 19 22 29 7 23 25 41 7 15 9 17 
14 1 4 5 6 18 19 22 29 7 23 25 41 27 28 
17 1 4 5 6 18 19 22 29 7 23 25 44 45 7 8 9 10 
10 1 4 5 6 36 37 34 35 20 21 
15 1 4 5 6 18 19 22 29 7 23 25 44 45 27 28 
17 1 4 5 6 18 19 22 29 7 23 25 18 19 7 8 9 10 
17 1 4 5 6 18 19 22 29 7 23 25 18 19 7 15 9 17 
15 1 4 5 6 18 19 22 29 7 23 25 18 19 27 28 
18 1 4 5 6 18 19 22 29 7 23 25 18 19 29 7 20 9 21 
17 1 4 5 6 18 19 22 29 7 23 25 30 31 7 8 9 10 
17 1 4 5 6 18 19 22 29 7 23 25 30 31 7 15 9 17 
15 1 4 5 6 18 19 22 29 7 23 25 30 31 27 28 
18 1 4 5 6 18 19 22 29 7 23 25 30 31 29 7 20 9 21 
17 1 4 5 6 18 19 22 29 7 23 25 46 47 7 8 9 10 
12 1 4 5 6 36 37 36 37 7 8 9 10 
15 1 4 5 6 18 19 22 29 7 23 25 46 47 27 28 
18 1 4 5 6 18 19 22 29 7 23 25 46 47 29 7 20 9 21 
20 1 4 5 6 18 19 22 29 7 23 25 22 29 7 23 25 7 8 9 10 
20 1 4 5 6 18 19 22 29 7 23 25 22 29 7 23 25 7 15 9 17 
18 1 4 5 6 18 19 22 29 7 23 25 22 29 7 23 25 27 28 
17 1 4 5 6 18 19 22 29 7 23 25 27 28 7 8 9 10 
17 1 4 5 6 18 19 22 29 7 23 25 27 28 7 15 9 17 
15 1 4 5 6 18 19 22 29 7 23 25 27 28 27 28 
17 1 4 5 6 18 19 22 29 7 23 25 13 32 7 8 9 10 
17 1 4 5 6 18 19 22 29 7 23 25 13 32 7 15 9 17 
10 1 4 5 6 44 45 7 8 9 10 
11 1 4 5 6 36 37 36 37 15 16 17 
15 1 4 5 6 18 19 22 29 7 23 25 13 32 27 28 
16 1 4 5 6 18 19 22 29 7 23 25 33 7 8 9 10 
14 1 4 5 6 18 19 22 29 7 23 25 33 27 28 
17 1 4 5 6 18 19 22 29 7 23 25 34 35 7 8 9 10 
16 1 4 5 6 18 19 22 29 7 23 25 34 35 15 16 17 
15 1 4 5 6 18 19 22 29 7 23 25 34 35 27 28 
15 1 4 5 6 18 19 22 29 7 23 25 34 35 20 21 
17 1 4 5 6 18 19 22 29 7 23 25 36 37 7 8 9 10 
16 1 4 5 6 18 19 22 29 7 23 25 36 37 15 16 17 
15 1 4 5 6 18 19 22 29 7 23 25 36 37 27 28 
10 1 4 5 6 36 37 36 37 27 28 
18 1 4 5 6 18 19 22 29 7 23 25 36 37 29 7 20 9 21 
17 1 4 5 6 18 19 22 29 7 23 25 38 39 7 8 9 10 
17 1 4 5 6 18 19 22 29 7 23 25 38 39 7 15 9 17 
15 1 4 5 6 18 19 22 29 7 23 25 38 39 27 28 
16 1 4 5 6 18 19 22 29 7 23 25 40 7 8 9 10 
14 1 4 5 6 18 19 22 29 7 23 25 40 27 28 
14 1 4 5 6 18 19 27 28 30 31 7 8 9 10 
14 1 4 5 6 18 19 27 28 30 31 7 15 9 17 
12 1 4 5 6 18 19 27 28 30 31 27 28 
15 1 4 5 6 18 19 27 28 30 31 29 7 20 9 21 
13 1 4 5 6 36 37 36 37 29 7 20 9 21 
14 1 4 5 6 18 19 27 28 27 28 7 8 9 10 
14 1 4 5 6 18 19 27 28 27 28 7 15 9 17 
12 1 4 5 6 18 19 27 28 27 28 27 28 
14 1 4 5 6 18 19 27 28 38 39 7 8 9 10 
14 1 4 5 6 18 19 27 28 38 39 7 15 9 17 
12 1 4 5 6 18 19 27 28 38 39 27 28 
14 1 4 5 6 18 19 13 32 42 43 7 8 9 10 
12 1 4 5 6 18 19 13 32 42 43 27 28 
13 1 4 5 6 18 19 13 32 41 7 8 9 10 
13 1 4 5 6 18 19 13 32 41 7 15 9 17 
12 1 4 5 6 36 37 38 39 7 8 9 10 
11 1 4 5 6 18 19 13 32 41 27 28 
14 1 4 5 6 18 19 13 32 44 45 7 8 9 10 
12 1 4 5 6 18 19 13 32 44 45 27 28 
14 1 4 5 6 18 19 13 32 30 31 7 8 9 10 
14 1 4 5 6 18 19 13 32 30 31 7 15 9 17 
12 1 4 5 6 18 19 13 32 30 31 27 28 
15 1 4 5 6 18 19 13 32 30 31 29 7 20 9 21 
14 1 4 5 6 18 19 13 32 46 47 7 8 9 10 
12 1 4 5 6 18 19 13 32 46 47 27 28 
15 1 4 5 6 18 19 13 32 46 47 29 7 20 9 21 
11 1 4 5 6 36 37 38 39 15 16 17 
14 1 4 5 6 18 19 13 32 27 28 7 8 9 10 
14 1 4 5 6 18 19 13 32 27 28 7 15 9 17 
12 1 4 5 6 18 19 13 32 27 28 27 28 
14 1 4 5 6 18 19 13 32 13 32 7 8 9 10 
14 1 4 5 6 18 19 13 32 13 32 7 15 9 17 
12 1 4 5 6 18 19 13 32 13 32 27 28 
13 1 4 5 6 18 19 13 32 33 7 8 9 10 
11 1 4 5 6 18 19 13 32 33 27 28 
14 1 4 5 6 18 19 13 32 36 37 7 8 9 10 
13 1 4 5 6 18 19 13 32 36 37 15 16 17 
10 1 4 5 6 36 37 38 39 27 28 
12 1 4 5 6 18 19 13 32 36 37 27 28 
15 1 4 5 6 18 19 13 32 36 37 29 7 20 9 21 
14 1 4 5 6 18 19 13 32 38 39 7 8 9 10 
14 1 4 5 6 18 19 13 32 38 39 7 15 9 17 
12 1 4 5 6 18 19 13 32 38 39 27 28 
13 1 4 5 6 18 19 13 32 40 7 8 9 10 
11 1 4 5 6 18 19 13 32 40 27 28 
13 1 4 5 6 18 19 33 42 43 7 8 9 10 
11 1 4 5 6 18 19 33 42 43 27 28 
13 1 4 5 6 18 19 33 44 45 7 8 9 10 
13 1 4 5 6 36 37 38 39 29 7 20 9 21 
11 1 4 5 6 18 19 33 44 45 27 28 
13 1 4 5 6 18 19 33 46 47 7 8 9 10 
11 1 4 5 6 18 19 33 46 47 27 28 
14 1 4 5 6 18 19 33 46 47 29 7 20 9 21 
13 1 4 5 6 18 19 33 27 28 7 8 9 10 
13 1 4 5 6 18 19 33 27 28 7 15 9 17 
11 1 4 5 6 18 19 33 27 28 27 28 
12 1 4 5 6 18 19 33 33 7 8 9 10 
10 1 4 5 6 18 19 33 33 27 28 
12 1 4 5 6 18 19 33 40 7 8 9 10 
11 1 4 5 6 36 37 40 7 8 9 10 
10 1 4 5 6 18 19 33 40 27 28 
14 1 4 5 6 18 19 36 37 42 43 7 8 9 10 
12 1 4 5 6 18 19 36 37 42 43 27 28 
16 1 4 5 6 18 19 36 37 11 12 13 14 7 8 9 10 
15 1 4 5 6 18 19 36 37 11 12 13 14 15 16 17 
14 1 4 5 6 18 19 36 37 11 12 13 14 27 28 
14 1 4 5 6 18 19 36 37 11 12 13 14 20 21 
13 1 4 5 6 18 19 36 37 41 7 8 9 10 
12 1 4 5 6 18 19 36 37 41 15 16 17 
11 1 4 5 6 18 19 36 37 41 27 28 
10 1 4 5 6 36 37 40 15 16 17 
14 1 4 5 6 18 19 36 37 44 45 7 8 9 10 
12 1 4 5 6 18 19 36 37 44 45 27 28 
14 1 4 5 6 18 19 36 37 30 31 7 8 9 10 
13 1 4 5 6 18 19 36 37 30 31 15 16 17 
12 1 4 5 6 18 19 36 37 30 31 27 28 
15 1 4 5 6 18 19 36 37 30 31 29 7 20 9 21 
14 1 4 5 6 18 19 36 37 46 47 7 8 9 10 
12 1 4 5 6 18 19 36 37 46 47 27 28 
12 1 4 5 6 18 19 36 37 46 47 20 21 
17 1 4 5 6 18 19 36 37 22 29 7 23 25 7 8 9 10 
9 1 4 5 6 36 37 40 27 28 
16 1 4 5 6 18 19 36 37 22 29 7 23 25 15 16 17 
15 1 4 5 6 18 19 36 37 22 29 7 23 25 27 28 
13 1 4 5 6 18 19 36 37 15 16 17 8 10 
14 1 4 5 6 18 19 36 37 15 16 17 15 16 17 
15 1 4 5 6 18 19 36 37 15 16 17 7 27 9 28 
16 1 4 5 6 18 19 36 37 15 16 17 29 7 20 9 21 
14 1 4 5 6 18 19 36 37 27 28 7 8 9 10 
13 1 4 5 6 18 19 36 37 27 28 15 16 17 
12 1 4 5 6 18 19 36 37 27 28 27 28 
13 1 4 5 6 18 19 36 37 33 7 8 9 10 
10 1 4 5 6 44 45 7 15 9 17 
12 1 4 5 6 36 37 40 29 7 20 9 21 
11 1 4 5 6 18 19 36 37 33 27 28 
14 1 4 5 6 18 19 36 37 34 35 7 8 9 10 
13 1 4 5 6 18 19 36 37 34 35 15 16 17 
12 1 4 5 6 18 19 36 37 34 35 27 28 
12 1 4 5 6 18 19 36 37 34 35 20 21 
14 1 4 5 6 18 19 36 37 36 37 7 8 9 10 
13 1 4 5 6 18 19 36 37 36 37 15 16 17 
12 1 4 5 6 18 19 36 37 36 37 27 28 
15 1 4 5 6 18 19 36 37 36 37 29 7 20 9 21 
14 1 4 5 6 18 19 36 37 38 39 7 8 9 10 
11 1 4 5 6 36 37 29 7 20 9 21 
13 1 4 5 6 18 19 36 37 38 39 15 16 17 
12 1 4 5 6 18 19 36 37 38 39 27 28 
13 1 4 5 6 18 19 36 37 40 7 8 9 10 
11 1 4 5 6 18 19 36 37 40 27 28 
14 1 4 5 6 18 19 38 39 42 43 7 8 9 10 
12 1 4 5 6 18 19 38 39 42 43 27 28 
14 1 4 5 6 18 19 38 39 44 45 7 8 9 10 
12 1 4 5 6 18 19 38 39 44 45 27 28 
14 1 4 5 6 18 19 38 39 30 31 7 8 9 10 
14 1 4 5 6 18 19 38 39 30 31 7 15 9 17 
11 1 4 5 6 36 37 29 7 20 9 21 
12 1 4 5 6 18 19 38 39 30 31 27 28 
15 1 4 5 6 18 19 38 39 30 31 29 7 20 9 21 
14 1 4 5 6 18 19 38 39 46 47 7 8 9 10 
12 1 4 5 6 18 19 38 39 46 47 27 28 
15 1 4 5 6 18 19 38 39 46 47 29 7 20 9 21 
17 1 4 5 6 18 19 38 39 22 29 7 23 25 7 8 9 10 
17 1 4 5 6 18 19 38 39 22 29 7 23 25 7 15 9 17 
15 1 4 5 6 18 19 38 39 22 29 7 23 25 27 28 
14 1 4 5 6 18 19 38 39 27 28 7 8 9 10 
14 1 4 5 6 18 19 38 39 27 28 7 15 9 17 
11 1 4 5 6 36 37 29 7 20 9 21 
12 1 4 5 6 18 19 38 39 27 28 27 28 
13 1 4 5 6 18 19 38 39 33 7 8 9 10 
11 1 4 5 6 18 19 38 39 33 27 28 
14 1 4 5 6 18 19 38 39 38 39 7 8 9 10 
14 1 4 5 6 18 19 38 39 38 39 7 15 9 17 
12 1 4 5 6 18 19 38 39 38 39 27 28 
13 1 4 5 6 18 19 38 39 40 7 8 9 10 
11 1 4 5 6 18 19 38 39 40 27 28 
13 1 4 5 6 18 19 40 42 43 7 8 9 10 
11 1 4 5 6 18 19 40 42 43 27 28 
11 1 4 5 6 36 37 29 7 20 9 21 
13 1 4 5 6 18 19 40 44 45 7 8 9 10 
11 1 4 5 6 18 19 40 44 45 27 28 
13 1 4 5 6 18 19 40 27 28 7 8 9 10 
13 1 4 5 6 18 19 40 27 28 7 15 9 17 
11 1 4 5 6 18 19 40 27 28 27 28 
12 1 4 5 6 18 19 40 40 7 8 9 10 
10 1 4 5 6 18 19 40 40 27 28 
14 1 4 5 6 30 31 42 43 42 43 7 8 9 10 
12 1 4 5 6 30 31 42 43 42 43 27 28 
16 1 4 5 6 30 31 42 43 11 12 13 14 7 8 9 10 
15 1 4 5 6 11 12 13 14 15 16 17 42 43 8 10 
15 1 4 5 6 30 31 42 43 11 12 13 14 15 16 17 
14 1 4 5 6 30 31 42 43 11 12 13 14 27 28 
14 1 4 5 6 30 31 42 43 11 12 13 14 20 21 
17 1 4 5 6 30 31 42 43 22 29 7 23 25 7 8 9 10 
17 1 4 5 6 30 31 42 43 22 29 7 23 25 7 15 9 17 
15 1 4 5 6 30 31 42 43 22 29 7 23 25 27 28 
14 1 4 5 6 30 31 42 43 27 28 7 8 9 10 
14 1 4 5 6 30 31 42 43 27 28 7 15 9 17 
12 1 4 5 6 30 31 42 43 27 28 27 28 
14 1 4 5 6 30 31 42 43 34 35 7 8 9 10 
16 1 4 5 6 11 12 13 14 15 16 17 42 43 15 16 17 
13 1 4 5 6 30 31 42 43 34 35 15 16 17 
12 1 4 5 6 30 31 42 43 34 35 27 28 
12 1 4 5 6 30 31 42 43 34 35 20 21 
14 1 4 5 6 30 31 44 45 42 43 7 8 9 10 
12 1 4 5 6 30 31 44 45 42 43 27 28 
16 1 4 5 6 30 31 44 45 11 12 13 14 7 8 9 10 
15 1 4 5 6 30 31 44 45 11 12 13 14 15 16 17 
14 1 4 5 6 30 31 44 45 11 12 13 14 27 28 
14 1 4 5 6 30 31 44 45 11 12 13 14 20 21 
14 1 4 5 6 30 31 44 45 44 45 7 8 9 10 
17 1 4 5 6 11 12 13 14 15 16 17 42 43 7 27 9 28 
12 1 4 5 6 30 31 44 45 44 45 27 28 
17 1 4 5 6 30 31 44 45 22 29 7 23 25 7 8 9 10 
17 1 4 5 6 30 31 44 45 22 29 7 23 25 7 15 9 17 
15 1 4 5 6 30 31 44 45 22 29 7 23 25 27 28 
14 1 4 5 6 30 31 44 45 27 28 7 8 9 10 
14 1 4 5 6 30 31 44 45 27 28 7 15 9 17 
12 1 4 5 6 30 31 44 45 27 28 27 28 
14 1 4 5 6 30 31 44 45 34 35 7 8 9 10 
13 1 4 5 6 30 31 44 45 34 35 15 16 17 
12 1 4 5 6 30 31 44 45 34 35 27 28 
18 1 4 5 6 11 12 13 14 15 16 17 42 43 29 7 20 9 21 
12 1 4 5 6 30 31 44 45 34 35 20 21 
14 1 4 5 6 30 31 30 31 42 43 7 8 9 10 
12 1 4 5 6 30 31 30 31 42 43 27 28 
14 1 4 5 6 30 31 30 31 44 45 7 8 9 10 
12 1 4 5 6 30 31 30 31 44 45 27 28 
14 1 4 5 6 30 31 30 31 30 31 7 8 9 10 
14 1 4 5 6 30 31 30 31 30 31 7 15 9 17 
12 1 4 5 6 30 31 30 31 30 31 27 28 
15 1 4 5 6 30 31 30 31 30 31 29 7 20 9 21 
14 1 4 5 6 30 31 30 31 46 47 7 8 9 10 
17 1 4 5 6 11 12 13 14 15 16 17 11 12 13 14 8 10 
12 1 4 5 6 30 31 30 31 46 47 27 28 
15 1 4 5 6 30 31 30 31 46 47 29 7 20 9 21 
17 1 4 5 6 30 31 30 31 22 29 7 23 25 7 8 9 10 
17 1 4 5 6 30 31 30 31 22 29 7 23 25 7 15 9 17 
15 1 4 5 6 30 31 30 31 22 29 7 23 25 27 28 
14 1 4 5 6 30 31 30 31 27 28 7 8 9 10 
14 1 4 5 6 30 31 30 31 27 28 7 15 9 17 
12 1 4 5 6 30 31 30 31 27 28 27 28 
13 1 4 5 6 30 31 30 31 33 7 8 9 10 
11 1 4 5 6 30 31 30 31 33 27 28 
8 1 4 5 6 44 45 27 28 
18 1 4 5 6 11 12 13 14 15 16 17 11 12 13 14 15 16 17 
13 1 4 5 6 30 31 30 31 40 7 8 9 10 
11 1 4 5 6 30 31 30 31 40 27 28 
14 1 4 5 6 30 31 46 47 42 43 7 8 9 10 
12 1 4 5 6 30 31 46 47 42 43 27 28 
16 1 4 5 6 30 31 46 47 11 12 13 14 7 8 9 10 
15 1 4 5 6 30 31 46 47 11 12 13 14 15 16 17 
14 1 4 5 6 30 31 46 47 11 12 13 14 27 28 
14 1 4 5 6 30 31 46 47 11 12 13 14 20 21 
14 1 4 5 6 30 31 46 47 44 45 7 8 9 10 
12 1 4 5 6 30 31 46 47 44 45 27 28 
19 1 4 5 6 11 12 13 14 15 16 17 11 12 13 14 7 27 9 28 
14 1 4 5 6 30 31 46 47 46 47 7 8 9 10 
12 1 4 5 6 30 31 46 47 46 47 27 28 
15 1 4 5 6 30 31 46 47 46 47 29 7 20 9 21 
17 1 4 5 6 30 31 46 47 22 29 7 23 25 7 8 9 10 
17 1 4 5 6 30 31 46 47 22 29 7 23 25 7 15 9 17 
15 1 4 5 6 30 31 46 47 22 29 7 23 25 27 28 
14 1 4 5 6 30 31 46 47 27 28 7 8 9 10 
14 1 4 5 6 30 31 46 47 27 28 7 15 9 17 
12 1 4 5 6 30 31 46 47 27 28 27 28 
14 1 4 5 6 30 31 46 47 34 35 7 8 9 10 
20 1 4 5 6 11 12 13 14 15 16 17 11 12 13 14 29 7 20 9 21 
13 1 4 5 6 30 31 46 47 34 35 15 16 17 
12 1 4 5 6 30 31 46 47 34 35 27 28 
12 1 4 5 6 30 31 46 47 34 35 20 21 
13 1 4 5 6 30 31 46 47 40 7 8 9 10 
11 1 4 5 6 30 31 46 47 40 27 28 
17 1 4 5 6 30 31 22 29 7 23 25 42 43 7 8 9 10 
15 1 4 5 6 30 31 22 29 7 23 25 42 43 27 28 
19 1 4 5 6 30 31 22 29 7 23 25 11 12 13 14 7 8 9 10 
18 1 4 5 6 30 31 22 29 7 23 25 11 12 13 14 15 16 17 
17 1 4 5 6 30 31 22 29 7 23 25 11 12 13 14 27 28 
15 1 4 5 6 11 12 13 14 15 16 17 8 10 8 10 
17 1 4 5 6 30 31 22 29 7 23 25 11 12 13 14 20 21 
16 1 4 5 6 30 31 22 29 7 23 25 41 7 8 9 10 
16 1 4 5 6 30 31 22 29 7 23 25 41 7 15 9 17 
14 1 4 5 6 30 31 22 29 7 23 25 41 27 28 
17 1 4 5 6 30 31 22 29 7 23 25 44 45 7 8 9 10 
15 1 4 5 6 30 31 22 29 7 23 25 44 45 27 28 
17 1 4 5 6 30 31 22 29 7 23 25 18 19 7 8 9 10 
17 1 4 5 6 30 31 22 29 7 23 25 18 19 7 15 9 17 
15 1 4 5 6 30 31 22 29 7 23 25 18 19 27 28 
18 1 4 5 6 30 31 22 29 7 23 25 18 19 29 7 20 9 21 
16 1 4 5 6 11 12 13 14 15 16 17 8 10 15 16 17 
17 1 4 5 6 30 31 22 29 7 23 25 30 31 7 8 9 10 
17 1 4 5 6 30 31 22 29 7 23 25 30 31 7 15 9 17 
15 1 4 5 6 30 31 22 29 7 23 25 30 31 27 28 
18 1 4 5 6 30 31 22 29 7 23 25 30 31 29 7 20 9 21 
17 1 4 5 6 30 31 22 29 7 23 25 46 47 7 8 9 10 
15 1 4 5 6 30 31 22 29 7 23 25 46 47 27 28 
18 1 4 5 6 30 31 22 29 7 23 25 46 47 29 7 20 9 21 
20 1 4 5 6 30 31 22 29 7 23 25 22 29 7 23 25 7 8 9 10 
20 1 4 5 6 30 31 22 29 7 23 25 22 29 7 23 25 7 15 9 17 
18 1 4 5 6 30 31 22 29 7 23 25 22 29 7 23 25 27 28 
17 1 4 5 6 11 12 13 14 15 16 17 8 10 7 27 9 28 
17 1 4 5 6 30 31 22 29 7 23 25 27 28 7 8 9 10 
17 1 4 5 6 30 31 22 29 7 23 25 27 28 7 15 9 17 
15 1 4 5 6 30 31 22 29 7 23 25 27 28 27 28 
17 1 4 5 6 30 31 22 29 7 23 25 13 32 7 8 9 10 
17 1 4 5 6 30 31 22 29 7 23 25 13 32 7 15 9 17 
15 1 4 5 6 30 31 22 29 7 23 25 13 32 27 28 
16 1 4 5 6 30 31 22 29 7 23 25 33 7 8 9 10 
14 1 4 5 6 30 31 22 29 7 23 25 33 27 28 
17 1 4 5 6 30 31 22 29 7 23 25 34 35 7 8 9 10 
16 1 4 5 6 30 31 22 29 7 23 25 34 35 15 16 17 
18 1 4 5 6 11 12 13 14 15 16 17 8 10 29 7 20 9 21 
15 1 4 5 6 30 31 22 29 7 23 25 34 35 27 28 
15 1 4 5 6 30 31 22 29 7 23 25 34 35 20 21 
17 1 4 5 6 30 31 22 29 7 23 25 36 37 7 8 9 10 
16 1 4 5 6 30 31 22 29 7 23 25 36 37 15 16 17 
15 1 4 5 6 30 31 22 29 7 23 25 36 37 27 28 
18 1 4 5 6 30 31 22 29 7 23 25 36 37 29 7 20 9 21 
17 1 4 5 6 30 31 22 29 7 23 25 38 39 7 8 9 10 
17 1 4 5 6 30 31 22 29 7 23 25 38 39 7 15 9 17 
15 1 4 5 6 30 31 22 29 7 23 25 38 39 27 28 
16 1 4 5 6 30 31 22 29 7 23 25 40 7 8 9 10 
14 1 4 5 6 11 12 13 14 15 16 17 41 8 10 
14 1 4 5 6 30 31 22 29 7 23 25 40 27 28 
14 1 4 5 6 30 31 27 28 30 31 7 8 9 10 
14 1 4 5 6 30 31 27 28 30 31 7 15 9 17 
12 1 4 5 6 30 31 27 28 30 31 27 28 
15 1 4 5 6 30 31 27 28 30 31 29 7 20 9 21 
14 1 4 5 6 30 31 27 28 27 28 7 8 9 10 
14 1 4 5 6 30 31 27 28 27 28 7 15 9 17 
12 1 4 5 6 30 31 27 28 27 28 27 28 
14 1 4 5 6 30 31 27 28 38 39 7 8 9 10 
14 1 4 5 6 30 31 27 28 38 39 7 15 9 17 
15 1 4 5 6 11 12 13 14 15 16 17 41 15 16 17 
12 1 4 5 6 30 31 27 28 38 39 27 28 
13 1 4 5 6 30 31 33 42 43 7 8 9 10 
11 1 4 5 6 30 31 33 42 43 27 28 
13 1 4 5 6 30 31 33 44 45 7 8 9 10 
11 1 4 5 6 30 31 33 44 45 27 28 
13 1 4 5 6 30 31 33 46 47 7 8 9 10 
11 1 4 5 6 30 31 33 46 47 27 28 
14 1 4 5 6 30 31 33 46 47 29 7 20 9 21 
13 1 4 5 6 30 31 33 27 28 7 8 9 10 
13 1 4 5 6 30 31 33 27 28 7 15 9 17 
16 1 4 5 6 11 12 13 14 15 16 17 41 7 27 9 28 
11 1 4 5 6 30 31 33 27 28 27 28 
12 1 4 5 6 30 31 33 33 7 8 9 10 
10 1 4 5 6 30 31 33 33 27 28 
12 1 4 5 6 30 31 33 40 7 8 9 10 
10 1 4 5 6 30 31 33 40 27 28 
13 1 4 5 6 30 31 40 42 43 7 8 9 10 
11 1 4 5 6 30 31 40 42 43 27 28 
13 1 4 5 6 30 31 40 44 45 7 8 9 10 
11 1 4 5 6 30 31 40 44 45 27 28 
13 1 4 5 6 30 31 40 27 28 7 8 9 10 
11 1 4 5 6 44 45 29 7 20 9 21 
17 1 4 5 6 11 12 13 14 15 16 17 41 29 7 20 9 21 
13 1 4 5 6 30 31 40 27 28 7 15 9 17 
11 1 4 5 6 30 31 40 27 28 27 28 
12 1 4 5 6 30 31 40 40 7 8 9 10 
10 1 4 5 6 30 31 40 40 27 28 
14 1 4 5 6 46 47 42 43 42 43 7 8 9 10 
12 1 4 5 6 46 47 42 43 42 43 27 28 
16 1 4 5 6 46 47 42 43 11 12 13 14 7 8 9 10 
15 1 4 5 6 46 47 42 43 11 12 13 14 15 16 17 
14 1 4 5 6 46 47 42 43 11 12 13 14 27 28 
14 1 4 5 6 46 47 42 43 11 12 13 14 20 21 
15 1 4 5 6 11 12 13 14 15 16 17 44 45 8 10 
17 1 4 5 6 46 47 42 43 22 29 7 23 25 7 8 9 10 
17 1 4 5 6 46 47 42 43 22 29 7 23 25 7 15 9 17 
15 1 4 5 6 46 47 42 43 22 29 7 23 25 27 28 
14 1 4 5 6 46 47 42 43 27 28 7 8 9 10 
14 1 4 5 6 46 47 42 43 27 28 7 15 9 17 
12 1 4 5 6 46 47 42 43 27 28 27 28 
14 1 4 5 6 46 47 42 43 34 35 7 8 9 10 
13 1 4 5 6 46 47 42 43 34 35 15 16 17 
12 1 4 5 6 46 47 42 43 34 35 27 28 
12 1 4 5 6 46 47 42 43 34 35 20 21 
16 1 4 5 6 11 12 13 14 15 16 17 44 45 15 16 17 
16 1 4 5 6 46 47 11 12 13 14 42 43 7 8 9 10 
14 1 4 5 6 46 47 11 12 13 14 42 43 27 28 
18 1 4 5 6 46 47 11 12 13 14 11 12 13 14 7 8 9 10 
17 1 4 5 6 46 47 11 12 13 14 11 12 13 14 15 16 17 
16 1 4 5 6 46 47 11 12 13 14 11 12 13 14 27 28 
16 1 4 5 6 46 47 11 12 13 14 11 12 13 14 20 21 
15 1 4 5 6 46 47 11 12 13 14 41 7 8 9 10 
14 1 4 5 6 46 47 11 12 13 14 41 15 16 17 
13 1 4 5 6 46 47 11 12 13 14 41 27 28 
16 1 4 5 6 46 47 11 12 13 14 44 45 7 8 9 10 
17 1 4 5 6 11 12 13 14 15 16 17 44 45 7 27 9 28 
14 1 4 5 6 46 47 11 12 13 14 44 45 27 28 
16 1 4 5 6 46 47 11 12 13 14 18 19 7 8 9 10 
15 1 4 5 6 46 47 11 12 13 14 18 19 15 16 17 
14 1 4 5 6 46 47 11 12 13 14 18 19 27 28 
14 1 4 5 6 46 47 11 12 13 14 18 19 20 21 
16 1 4 5 6 46 47 11 12 13 14 30 31 7 8 9 10 
15 1 4 5 6 46 47 11 12 13 14 30 31 15 16 17 
14 1 4 5 6 46 47 11 12 13 14 30 31 27 28 
14 1 4 5 6 46 47 11 12 13 14 30 31 20 21 
16 1 4 5 6 46 47 11 12 13 14 46 47 7 8 9 10 
18 1 4 5 6 11 12 13 14 15 16 17 44 45 29 7 20 9 21 
14 1 4 5 6 46 47 11 12 13 14 46 47 27 28 
14 1 4 5 6 46 47 11 12 13 14 46 47 20 21 
19 1 4 5 6 46 47 11 12 13 14 22 23 26 24 25 7 8 9 10 
18 1 4 5 6 46 47 11 12 13 14 22 23 24 25 7 8 9 10 
18 1 4 5 6 46 47 11 12 13 14 22 23 26 24 25 15 16 17 
17 1 4 5 6 46 47 11 12 13 14 22 23 24 25 15 16 17 
17 1 4 5 6 46 47 11 12 13 14 22 23 26 24 25 27 28 
16 1 4 5 6 46 47 11 12 13 14 22 23 24 25 27 28 
15 1 4 5 6 46 47 11 12 13 14 15 16 17 8 10 
16 1 4 5 6 46 47 11 12 13 14 15 16 17 15 16 17 
17 1 4 5 6 11 12 13 14 15 16 17 18 19 7 8 9 10 
17 1 4 5 6 46 47 11 12 13 14 15 16 17 7 27 9 28 
18 1 4 5 6 46 47 11 12 13 14 15 16 17 29 7 20 9 21 
16 1 4 5 6 46 47 11 12 13 14 27 28 7 8 9 10 
15 1 4 5 6 46 47 11 12 13 14 27 28 15 16 17 
14 1 4 5 6 46 47 11 12 13 14 27 28 27 28 
16 1 4 5 6 46 47 11 12 13 14 13 32 7 8 9 10 
15 1 4 5 6 46 47 11 12 13 14 13 32 15 16 17 
14 1 4 5 6 46 47 11 12 13 14 13 32 27 28 
15 1 4 5 6 46 47 11 12 13 14 33 7 8 9 10 
13 1 4 5 6 46 47 11 12 13 14 33 27 28 
16 1 4 5 6 11 12 13 14 15 16 17 18 19 15 16 17 
16 1 4 5 6 46 47 11 12 13 14 34 35 7 8 9 10 
15 1 4 5 6 46 47 11 12 13 14 34 35 15 16 17 
14 1 4 5 6 46 47 11 12 13 14 34 35 27 28 
14 1 4 5 6 46 47 11 12 13 14 34 35 20 21 
16 1 4 5 6 46 47 11 12 13 14 36 37 7 8 9 10 
15 1 4 5 6 46 47 11 12 13 14 36 37 15 16 17 
14 1 4 5 6 46 47 11 12 13 14 36 37 27 28 
14 1 4 5 6 46 47 11 12 13 14 36 37 20 21 
16 1 4 5 6 46 47 11 12 13 14 38 39 7 8 9 10 
15 1 4 5 6 46 47 11 12 13 14 38 39 15 16 17 
17 1 4 5 6 11 12 13 14 15 16 17 18 19 7 27 9 28 
14 1 4 5 6 46 47 11 12 13 14 38 39 27 28 
15 1 4 5 6 46 47 11 12 13 14 40 7 8 9 10 
13 1 4 5 6 46 47 11 12 13 14 40 27 28 
16 1 4 5 6 46 47 11 12 13 14 20 21 7 8 9 10 
15 1 4 5 6 46 47 11 12 13 14 20 21 15 16 17 
14 1 4 5 6 46 47 11 12 13 14 20 21 27 28 
14 1 4 5 6 46 47 11 12 13 14 20 21 20 21 
14 1 4 5 6 46 47 44 45 42 43 7 8 9 10 
12 1 4 5 6 46 47 44 45 42 43 27 28 
16 1 4 5 6 46 47 44 45 11 12 13 14 7 8 9 10 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 29 7 20 9 21 
15 1 4 5 6 46 47 44 45 11 12 13 14 15 16 17 
14 1 4 5 6 46 47 44 45 11 12 13 14 27 28 
14 1 4 5 6 46 47 44 45 11 12 13 14 20 21 
14 1 4 5 6 46 47 44 45 44 45 7 8 9 10 
12 1 4 5 6 46 47 44 45 44 45 27 28 
17 1 4 5 6 46 47 44 45 22 29 7 23 25 7 8 9 10 
17 1 4 5 6 46 47 44 45 22 29 7 23 25 7 15 9 17 
15 1 4 5 6 46 47 44 45 22 29 7 23 25 27 28 
14 1 4 5 6 46 47 44 45 27 28 7 8 9 10 
14 1 4 5 6 46 47 44 45 27 28 7 15 9 17 
15 1 4 5 6 11 12 13 14 15 16 17 30 31 8 10 
12 1 4 5 6 46 47 44 45 27 28 27 28 
14 1 4 5 6 46 47 44 45 34 35 7 8 9 10 
13 1 4 5 6 46 47 44 45 34 35 15 16 17 
12 1 4 5 6 46 47 44 45 34 35 27 28 
12 1 4 5 6 46 47 44 45 34 35 20 21 
14 1 4 5 6 46 47 46 47 42 43 7 8 9 10 
12 1 4 5 6 46 47 46 47 42 43 27 28 
16 1 4 5 6 46 47 46 47 11 12 13 14 7 8 9 10 
15 1 4 5 6 46 47 46 47 11 12 13 14 15 16 17 
14 1 4 5 6 46 47 46 47 11 12 13 14 27 28 
10 1 4 5 6 18 19 7 8 9 10 
16 1 4 5 6 11 12 13 14 15 16 17 30 31 15 16 17 
14 1 4 5 6 46 47 46 47 11 12 13 14 20 21 
14 1 4 5 6 46 47 46 47 44 45 7 8 9 10 
12 1 4 5 6 46 47 46 47 44 45 27 28 
14 1 4 5 6 46 47 46 47 46 47 7 8 9 10 
12 1 4 5 6 46 47 46 47 46 47 27 28 
15 1 4 5 6 46 47 46 47 46 47 29 7 20 9 21 
17 1 4 5 6 46 47 46 47 22 29 7 23 25 7 8 9 10 
17 1 4 5 6 46 47 46 47 22 29 7 23 25 7 15 9 17 
15 1 4 5 6 46 47 46 47 22 29 7 23 25 27 28 
14 1 4 5 6 46 47 46 47 27 28 7 8 9 10 
17 1 4 5 6 11 12 13 14 15 16 17 30 31 7 27 9 28 
14 1 4 5 6 46 47 46 47 27 28 7 15 9 17 
12 1 4 5 6 46 47 46 47 27 28 27 28 
14 1 4 5 6 46 47 46 47 34 35 7 8 9 10 
13 1 4 5 6 46 47 46 47 34 35 15 16 17 
12 1 4 5 6 46 47 46 47 34 35 27 28 
12 1 4 5 6 46 47 46 47 34 35 20 21 
13 1 4 5 6 46 47 46 47 40 7 8 9 10 
11 1 4 5 6 46 47 46 47 40 27 28 
17 1 4 5 6 46 47 22 29 7 23 25 42 43 7 8 9 10 
15 1 4 5 6 46 47 22 29 7 23 25 42 43 27 28 
18 1 4 5 6 11 12 13 14 15 16 17 30 31 29 7 20 9 21 
19 1 4 5 6 46 47 22 29 7 23 25 11 12 13 14 7 8 9 10 
18 1 4 5 6 46 47 22 29 7 23 25 11 12 13 14 15 16 17 
17 1 4 5 6 46 47 22 29 7 23 25 11 12 13 14 27 28 
17 1 4 5 6 46 47 22 29 7 23 25 11 12 13 14 20 21 
16 1 4 5 6 46 47 22 29 7 23 25 41 7 8 9 10 
16 1 4 5 6 46 47 22 29 7 23 25 41 7 15 9 17 
14 1 4 5 6 46 47 22 29 7 23 25 41 27 28 
17 1 4 5 6 46 47 22 29 7 23 25 44 45 7 8 9 10 
15 1 4 5 6 46 47 22 29 7 23 25 44 45 27 28 
17 1 4 5 6 46 47 22 29 7 23 25 18 19 7 8 9 10 
15 1 4 5 6 11 12 13 14 15 16 17 46 47 8 10 
17 1 4 5 6 46 47 22 29 7 23 25 18 19 7 15 9 17 
15 1 4 5 6 46 47 22 29 7 23 25 18 19 27 28 
18 1 4 5 6 46 47 22 29 7 23 25 18 19 29 7 20 9 21 
17 1 4 5 6 46 47 22 29 7 23 25 30 31 7 8 9 10 
17 1 4 5 6 46 47 22 29 7 23 25 30 31 7 15 9 17 
15 1 4 5 6 46 47 22 29 7 23 25 30 31 27 28 
18 1 4 5 6 46 47 22 29 7 23 25 30 31 29 7 20 9 21 
17 1 4 5 6 46 47 22 29 7 23 25 46 47 7 8 9 10 
15 1 4 5 6 46 47 22 29 7 23 25 46 47 27 28 
18 1 4 5 6 46 47 22 29 7 23 25 46 47 29 7 20 9 21 
16 1 4 5 6 11 12 13 14 15 16 17 46 47 15 16 17 
20 1 4 5 6 46 47 22 29 7 23 25 22 29 7 23 25 7 8 9 10 
20 1 4 5 6 46 47 22 29 7 23 25 22 29 7 23 25 7 15 9 17 
18 1 4 5 6 46 47 22 29 7 23 25 22 29 7 23 25 27 28 
17 1 4 5 6 46 47 22 29 7 23 25 27 28 7 8 9 10 
17 1 4 5 6 46 47 22 29 7 23 25 27 28 7 15 9 17 
15 1 4 5 6 46 47 22 29 7 23 25 27 28 27 28 
17 1 4 5 6 46 47 22 29 7 23 25 13 32 7 8 9 10 
17 1 4 5 6 46 47 22 29 7 23 25 13 32 7 15 9 17 
15 1 4 5 6 46 47 22 29 7 23 25 13 32 27 28 
16 1 4 5 6 46 47 22 29 7 23 25 33 7 8 9 10 
17 1 4 5 6 11 12 13 14 15 16 17 46 47 7 27 9 28 
14 1 4 5 6 46 47 22 29 7 23 25 33 27 28 
17 1 4 5 6 46 47 22 29 7 23 25 34 35 7 8 9 10 
16 1 4 5 6 46 47 22 29 7 23 25 34 35 15 16 17 
15 1 4 5 6 46 47 22 29 7 23 25 34 35 27 28 
15 1 4 5 6 46 47 22 29 7 23 25 34 35 20 21 
17 1 4 5 6 46 47 22 29 7 23 25 36 37 7 8 9 10 
16 1 4 5 6 46 47 22 29 7 23 25 36 37 15 16 17 
15 1 4 5 6 46 47 22 29 7 23 25 36 37 27 28 
15 1 4 5 6 46 47 22 29 7 23 25 36 37 20 21 
18 1 4 5 6 36 37 22 29 7 23 25 36 37 29 7 20 9 21 
18 1 4 5 6 11 12 13 14 15 16 17 46 47 29 7 20 9 21 
23 1 4 5 6 11 12 13 14 15 16 17 22 29 7 23 25 36 37 29 7 20 9 21 
25 1 4 5 6 11 12 13 14 15 16 17 18 19 22 29 7 23 25 36 37 29 7 20 9 21 
24 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 22 29 7 23 25 36 37 20 21 
9 1 4 5 6 29 7 20 9 21 
8 1 4 5 6 7 8 9 10 
17 1 4 5 6 41 22 29 7 23 25 36 37 29 7 20 9 21 
21 1 4 5 6 22 29 7 23 25 22 29 7 23 25 36 37 29 7 20 9 21 
18 1 4 5 6 11 12 13 14 15 16 17 22 29 7 23 25 8 10 
19 1 4 5 6 11 12 13 14 15 16 17 22 29 7 23 25 15 16 17 
20 1 4 5 6 11 12 13 14 15 16 17 22 29 7 23 25 7 27 9 28 
10 1 4 5 6 18 19 7 15 9 17 
21 1 4 5 6 11 12 13 14 15 16 17 22 29 7 23 25 29 7 20 9 21 
16 1 4 5 6 11 12 13 14 15 16 17 15 16 17 8 10 
17 1 4 5 6 11 12 13 14 15 16 17 15 16 17 15 16 17 
18 1 4 5 6 11 12 13 14 15 16 17 15 16 17 7 27 9 28 
19 1 4 5 6 11 12 13 14 15 16 17 15 16 17 29 7 20 9 21 
15 1 4 5 6 11 12 13 14 15 16 17 7 27 9 28 
15 1 4 5 6 11 12 13 14 15 16 17 7 27 9 28 
15 1 4 5 6 11 12 13 14 15 16 17 7 27 9 28 
15 1 4 5 6 11 12 13 14 15 16 17 7 27 9 28 
15 1 4 5 6 11 12 13 14 15 16 17 13 32 8 10 
8 1 4 5 6 18 19 27 28 
16 1 4 5 6 11 12 13 14 15 16 17 13 32 15 16 17 
17 1 4 5 6 11 12 13 14 15 16 17 13 32 7 27 9 28 
18 1 4 5 6 11 12 13 14 15 16 17 13 32 29 7 20 9 21 
14 1 4 5 6 11 12 13 14 15 16 17 33 8 10 
15 1 4 5 6 11 12 13 14 15 16 17 33 15 16 17 
16 1 4 5 6 11 12 13 14 15 16 17 33 7 27 9 28 
17 1 4 5 6 11 12 13 14 15 16 17 33 29 7 20 9 21 
15 1 4 5 6 11 12 13 14 15 16 17 34 35 8 10 
16 1 4 5 6 11 12 13 14 15 16 17 34 35 15 16 17 
17 1 4 5 6 11 12 13 14 15 16 17 34 35 7 27 9 28 
11 1 4 5 6 18 19 29 7 20 9 21 
18 1 4 5 6 11 12 13 14 15 16 17 34 35 29 7 20 9 21 
15 1 4 5 6 11 12 13 14 15 16 17 36 37 8 10 
16 1 4 5 6 11 12 13 14 15 16 17 36 37 15 16 17 
17 1 4 5 6 11 12 13 14 15 16 17 36 37 7 27 9 28 
18 1 4 5 6 11 12 13 14 15 16 17 36 37 29 7 20 9 21 
15 1 4 5 6 11 12 13 14 15 16 17 38 39 8 10 
16 1 4 5 6 11 12 13 14 15 16 17 38 39 15 16 17 
17 1 4 5 6 11 12 13 14 15 16 17 38 39 7 27 9 28 
18 1 4 5 6 11 12 13 14 15 16 17 38 39 29 7 20 9 21 
14 1 4 5 6 11 12 13 14 15 16 17 40 8 10 
10 1 4 5 6 30 31 7 8 9 10 
15 1 4 5 6 11 12 13 14 15 16 17 40 15 16 17 
16 1 4 5 6 11 12 13 14 15 16 17 40 7 27 9 28 
17 1 4 5 6 11 12 13 14 15 16 17 40 29 7 20 9 21 
16 1 4 5 6 11 12 13 14 15 16 17 29 7 20 9 21 
16 1 4 5 6 11 12 13 14 15 16 17 29 7 20 9 21 
16 1 4 5 6 11 12 13 14 15 16 17 29 7 20 9 21 
16 1 4 5 6 11 12 13 14 15 16 17 29 7 20 9 21 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 42 43 7 8 9 10 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 42 43 15 16 17 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 42 43 7 27 9 28 
6 1 4 5 6 27 28 
10 1 4 5 6 30 31 7 15 9 17 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 42 43 29 7 20 9 21 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 11 12 13 14 7 8 9 10 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 11 12 13 14 15 16 17 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 11 12 13 14 7 27 9 28 
22 1 4 5 6 11 12 13 14 15 16 17 18 19 11 12 13 14 29 7 20 9 21 
17 1 4 5 6 11 12 13 14 15 16 17 18 19 7 8 9 10 
17 1 4 5 6 11 12 13 14 15 16 17 18 19 7 8 9 10 
17 1 4 5 6 11 12 13 14 15 16 17 18 19 7 8 9 10 
17 1 4 5 6 11 12 13 14 15 16 17 18 19 7 8 9 10 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 41 7 8 9 10 
8 1 4 5 6 30 31 27 28 
17 1 4 5 6 11 12 13 14 15 16 17 18 19 41 15 16 17 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 41 7 27 9 28 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 41 29 7 20 9 21 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 44 45 7 8 9 10 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 44 45 15 16 17 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 44 45 7 27 9 28 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 44 45 29 7 20 9 21 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 18 19 7 8 9 10 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 18 19 15 16 17 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 18 19 7 27 9 28 
11 1 4 5 6 30 31 29 7 20 9 21 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 18 19 29 7 20 9 21 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 7 8 9 10 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 15 16 17 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 7 27 9 28 
17 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 20 21 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 46 47 7 8 9 10 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 46 47 15 16 17 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 46 47 7 27 9 28 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 46 47 29 7 20 9 21 
22 1 4 5 6 11 12 13 14 15 16 17 18 19 22 29 7 23 25 7 8 9 10 
10 1 4 5 6 46 47 7 8 9 10 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 22 29 7 23 25 15 16 17 
22 1 4 5 6 11 12 13 14 15 16 17 18 19 22 29 7 23 25 7 27 9 28 
23 1 4 5 6 11 12 13 14 15 16 17 18 19 22 29 7 23 25 29 7 20 9 21 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 15 16 17 8 10 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 15 16 17 15 16 17 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 15 16 17 7 27 9 28 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 15 16 17 29 7 20 9 21 
17 1 4 5 6 11 12 13 14 15 16 17 18 19 7 27 9 28 
17 1 4 5 6 11 12 13 14 15 16 17 18 19 7 27 9 28 
17 1 4 5 6 11 12 13 14 15 16 17 18 19 7 27 9 28 
10 1 4 5 6 46 47 7 15 9 17 
17 1 4 5 6 11 12 13 14 15 16 17 18 19 7 27 9 28 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 13 32 7 8 9 10 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 13 32 15 16 17 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 13 32 7 27 9 28 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 13 32 29 7 20 9 21 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 33 7 8 9 10 
17 1 4 5 6 11 12 13 14 15 16 17 18 19 33 15 16 17 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 33 7 27 9 28 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 33 29 7 20 9 21 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 34 35 7 8 9 10 
8 1 4 5 6 46 47 27 28 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 34 35 15 16 17 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 34 35 7 27 9 28 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 34 35 29 7 20 9 21 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 36 37 7 8 9 10 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 36 37 15 16 17 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 36 37 7 27 9 28 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 36 37 29 7 20 9 21 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 38 39 7 8 9 10 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 38 39 15 16 17 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 38 39 7 27 9 28 
11 1 4 5 6 46 47 29 7 20 9 21 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 38 39 29 7 20 9 21 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 40 7 8 9 10 
17 1 4 5 6 11 12 13 14 15 16 17 18 19 40 15 16 17 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 40 7 27 9 28 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 40 29 7 20 9 21 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 29 7 20 9 21 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 29 7 20 9 21 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 29 7 20 9 21 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 29 7 20 9 21 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 42 43 7 8 9 10 
13 1 4 5 6 22 29 7 23 25 7 8 9 10 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 42 43 15 16 17 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 42 43 7 27 9 28 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 42 43 20 21 
23 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 11 12 13 14 7 8 9 10 
22 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 11 12 13 14 15 16 17 
23 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 11 12 13 14 7 27 9 28 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 11 12 13 14 20 21 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 7 8 9 10 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 7 8 9 10 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 7 8 9 10 
13 1 4 5 6 22 29 7 23 25 7 15 9 17 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 7 8 9 10 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 41 7 8 9 10 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 41 15 16 17 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 41 7 27 9 28 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 41 20 21 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 44 45 7 8 9 10 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 44 45 15 16 17 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 44 45 7 27 9 28 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 44 45 20 21 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 18 19 7 8 9 10 
11 1 4 5 6 22 29 7 23 25 27 28 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 18 19 15 16 17 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 18 19 7 27 9 28 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 18 19 20 21 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 30 31 7 8 9 10 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 30 31 15 16 17 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 30 31 7 27 9 28 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 30 31 20 21 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 46 47 7 8 9 10 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 46 47 15 16 17 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 46 47 7 27 9 28 
9 1 4 5 6 29 7 20 9 21 
14 1 4 5 6 22 29 7 23 25 29 7 20 9 21 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 46 47 20 21 
24 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 22 29 7 23 25 7 8 9 10 
23 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 22 29 7 23 25 15 16 17 
24 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 22 29 7 23 25 7 27 9 28 
22 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 22 29 7 23 25 20 21 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 15 16 17 8 10 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 15 16 17 15 16 17 
22 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 15 16 17 7 27 9 28 
23 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 15 16 17 29 7 20 9 21 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 7 27 9 28 
8 1 4 5 6 7 15 9 17 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 7 27 9 28 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 7 27 9 28 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 7 27 9 28 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 13 32 7 8 9 10 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 13 32 15 16 17 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 13 32 7 27 9 28 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 13 32 20 21 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 33 7 8 9 10 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 33 15 16 17 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 33 7 27 9 28 
8 1 4 5 6 7 15 9 17 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 33 20 21 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 34 35 7 8 9 10 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 34 35 15 16 17 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 34 35 7 27 9 28 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 34 35 20 21 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 36 37 7 8 9 10 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 36 37 15 16 17 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 36 37 7 27 9 28 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 36 37 20 21 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 38 39 7 8 9 10 
8 1 4 5 6 7 15 9 17 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 38 39 15 16 17 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 38 39 27 28 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 38 39 20 21 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 40 7 8 9 10 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 40 15 16 17 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 40 7 27 9 28 
18 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 40 20 21 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 20 21 7 8 9 10 
20 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 20 21 15 16 17 
21 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 20 21 7 27 9 28 
8 1 4 5 6 7 15 9 17 
19 1 4 5 6 11 12 13 14 15 16 17 18 19 30 31 20 21 20 21 
12 1 4 5 6 42 43 42 43 7 8 9 10 
10 1 4 5 6 42 43 42 43 27 28 
14 1 4 5 6 42 43 11 12 13 14 7 8 9 10 
13 1 4 5 6 42 43 11 12 13 14 15 16 17 
12 1 4 5 6 42 43 11 12 13 14 27 28 
12 1 4 5 6 42 43 11 12 13 14 20 21 
15 1 4 5 6 42 43 22 29 7 23 25 7 8 9 10 
15 1 4 5 6 42 43 22 29 7 23 25 7 15 9 17 
13 1 4 5 6 42 43 22 29 7 23 25 27 28 
10 1 4 5 6 27 28 7 8 9 10 
12 1 4 5 6 42 43 27 28 7 8 9 10 
12 1 4 5 6 42 43 27 28 7 15 9 17 
10 1 4 5 6 42 43 27 28 27 28 
12 1 4 5 6 42 43 34 35 7 8 9 10 
11 1 4 5 6 42 43 34 35 15 16 17 
10 1 4 5 6 42 43 34 35 27 28 
10 1 4 5 6 42 43 34 35 20 21 
11 1 4 5 6 41 42 43 7 8 9 10 
9 1 4 5 6 41 42 43 27 28 
10 1 4 5 6 41 41 7 8 9 10 
10 1 4 5 6 27 28 7 15 9 17 
10 1 4 5 6 41 41 7 15 9 17 
8 1 4 5 6 41 41 27 28 
11 1 4 5 6 41 44 45 7 8 9 10 
9 1 4 5 6 41 44 45 27 28 
11 1 4 5 6 41 30 31 7 8 9 10 
11 1 4 5 6 41 30 31 7 15 9 17 
9 1 4 5 6 41 30 31 27 28 
12 1 4 5 6 41 30 31 29 7 20 9 21 
11 1 4 5 6 41 46 47 7 8 9 10 
9 1 4 5 6 41 46 47 27 28 
8 1 4 5 6 27 28 27 28 
12 1 4 5 6 41 46 47 29 7 20 9 21 
11 1 4 5 6 41 27 28 7 8 9 10 
11 1 4 5 6 41 27 28 7 15 9 17 
9 1 4 5 6 41 27 28 27 28 
10 1 4 5 6 41 33 7 8 9 10 
8 1 4 5 6 41 33 27 28 
11 1 4 5 6 41 38 39 7 8 9 10 
11 1 4 5 6 41 38 39 7 15 9 17 
9 1 4 5 6 41 38 39 27 28 
10 1 4 5 6 41 40 7 8 9 10 
11 1 4 5 6 27 28 29 7 20 9 21 
8 1 4 5 6 41 40 27 28 
12 1 4 5 6 44 45 42 43 7 8 9 10 
10 1 4 5 6 44 45 42 43 27 28 
14 1 4 5 6 44 45 11 12 13 14 7 8 9 10 
13 1 4 5 6 44 45 11 12 13 14 15 16 17 
12 1 4 5 6 44 45 11 12 13 14 27 28 
12 1 4 5 6 44 45 11 12 13 14 20 21 
12 1 4 5 6 44 45 44 45 7 8 9 10 
10 1 4 5 6 44 45 44 45 27 28 
15 1 4 5 6 44 45 22 29 7 23 25 7 8 9 10 
10 1 4 5 6 13 32 7 8 9 10 
15 1 4 5 6 44 45 22 29 7 23 25 7 15 9 17 
13 1 4 5 6 44 45 22 29 7 23 25 27 28 
12 1 4 5 6 44 45 27 28 7 8 9 10 
12 1 4 5 6 44 45 27 28 7 15 9 17 
10 1 4 5 6 44 45 27 28 27 28 
12 1 4 5 6 44 45 34 35 7 8 9 10 
11 1 4 5 6 44 45 34 35 15 16 17 
10 1 4 5 6 44 45 34 35 27 28 
10 1 4 5 6 44 45 34 35 20 21 
12 1 4 5 6 18 19 42 43 7 8 9 10 
10 1 4 5 6 42 43 7 8 9 10 
10 1 4 5 6 13 32 7 15 9 17 
10 1 4 5 6 18 19 42 43 27 28 
11 1 4 5 6 18 19 41 7 8 9 10 
11 1 4 5 6 18 19 41 7 15 9 17 
9 1 4 5 6 18 19 41 27 28 
12 1 4 5 6 18 19 44 45 7 8 9 10 
10 1 4 5 6 18 19 44 45 27 28 
12 1 4 5 6 18 19 18 19 7 8 9 10 
12 1 4 5 6 18 19 18 19 7 15 9 17 
10 1 4 5 6 18 19 18 19 27 28 
13 1 4 5 6 18 19 18 19 29 7 20 9 21 
8 1 4 5 6 13 32 27 28 
12 1 4 5 6 18 19 30 31 7 8 9 10 
12 1 4 5 6 18 19 30 31 7 15 9 17 
10 1 4 5 6 18 19 30 31 27 28 
13 1 4 5 6 18 19 30 31 29 7 20 9 21 
12 1 4 5 6 18 19 46 47 7 8 9 10 
10 1 4 5 6 18 19 46 47 27 28 
13 1 4 5 6 18 19 46 47 29 7 20 9 21 
15 1 4 5 6 18 19 22 29 7 23 25 7 8 9 10 
15 1 4 5 6 18 19 22 29 7 23 25 7 15 9 17 
13 1 4 5 6 18 19 22 29 7 23 25 27 28 
11 1 4 5 6 13 32 29 7 20 9 21 
12 1 4 5 6 18 19 27 28 7 8 9 10 
12 1 4 5 6 18 19 27 28 7 15 9 17 
10 1 4 5 6 18 19 27 28 27 28 
12 1 4 5 6 18 19 13 32 7 8 9 10 
12 1 4 5 6 18 19 13 32 7 15 9 17 
10 1 4 5 6 18 19 13 32 27 28 
11 1 4 5 6 18 19 33 7 8 9 10 
9 1 4 5 6 18 19 33 27 28 
12 1 4 5 6 18 19 36 37 7 8 9 10 
11 1 4 5 6 18 19 36 37 15 16 17 
9 1 4 5 6 33 7 8 9 10 
10 1 4 5 6 18 19 36 37 27 28 
13 1 4 5 6 18 19 36 37 29 7 20 9 21 
12 1 4 5 6 18 19 38 39 7 8 9 10 
12 1 4 5 6 18 19 38 39 7 15 9 17 
10 1 4 5 6 18 19 38 39 27 28 
11 1 4 5 6 18 19 40 7 8 9 10 
9 1 4 5 6 18 19 40 27 28 
12 1 4 5 6 30 31 42 43 7 8 9 10 
10 1 4 5 6 30 31 42 43 27 28 
12 1 4 5 6 30 31 44 45 7 8 9 10 
9 1 4 5 6 33 7 15 9 17 
10 1 4 5 6 30 31 44 45 27 28 
12 1 4 5 6 30 31 30 31 7 8 9 10 
12 1 4 5 6 30 31 30 31 7 15 9 17 
10 1 4 5 6 30 31 30 31 27 28 
13 1 4 5 6 30 31 30 31 29 7 20 9 21 
12 1 4 5 6 30 31 46 47 7 8 9 10 
10 1 4 5 6 30 31 46 47 27 28 
13 1 4 5 6 30 31 46 47 29 7 20 9 21 
15 1 4 5 6 30 31 22 29 7 23 25 7 8 9 10 
15 1 4 5 6 30 31 22 29 7 23 25 7 15 9 17 
7 1 4 5 6 33 27 28 
13 1 4 5 6 30 31 22 29 7 23 25 27 28 
12 1 4 5 6 30 31 27 28 7 8 9 10 
12 1 4 5 6 30 31 27 28 7 15 9 17 
10 1 4 5 6 30 31 27 28 27 28 
11 1 4 5 6 30 31 33 7 8 9 10 
9 1 4 5 6 30 31 33 27 28 
11 1 4 5 6 30 31 40 7 8 9 10 
9 1 4 5 6 30 31 40 27 28 
12 1 4 5 6 46 47 42 43 7 8 9 10 
10 1 4 5 6 46 47 42 43 27 28 
10 1 4 5 6 33 29 7 20 9 21 
14 1 4 5 6 46 47 11 12 13 14 7 8 9 10 
13 1 4 5 6 46 47 11 12 13 14 15 16 17 
12 1 4 5 6 46 47 11 12 13 14 27 28 
12 1 4 5 6 46 47 11 12 13 14 20 21 
12 1 4 5 6 46 47 44 45 7 8 9 10 
10 1 4 5 6 46 47 44 45 27 28 
12 1 4 5 6 46 47 46 47 7 8 9 10 
10 1 4 5 6 46 47 46 47 27 28 
13 1 4 5 6 46 47 46 47 29 7 20 9 21 
15 1 4 5 6 46 47 22 29 7 23 25 7 8 9 10 
10 1 4 5 6 34 35 7 8 9 10 
15 1 4 5 6 46 47 22 29 7 23 25 7 15 9 17 
13 1 4 5 6 46 47 22 29 7 23 25 27 28 
12 1 4 5 6 46 47 27 28 7 8 9 10 
12 1 4 5 6 46 47 27 28 7 15 9 17 
10 1 4 5 6 46 47 27 28 27 28 
12 1 4 5 6 46 47 34 35 7 8 9 10 
11 1 4 5 6 46 47 34 35 15 16 17 
10 1 4 5 6 46 47 34 35 27 28 
10 1 4 5 6 46 47 34 35 20 21 
11 1 4 5 6 46 47 40 7 8 9 10 
9 1 4 5 6 34 35 15 16 17 
9 1 4 5 6 46 47 40 27 28 
15 1 4 5 6 22 29 7 23 25 42 43 7 8 9 10 
13 1 4 5 6 22 29 7 23 25 42 43 27 28 
17 1 4 5 6 22 29 7 23 25 11 12 13 14 7 8 9 10 
16 1 4 5 6 22 29 7 23 25 11 12 13 14 15 16 17 
15 1 4 5 6 22 29 7 23 25 11 12 13 14 27 28 
15 1 4 5 6 22 29 7 23 25 11 12 13 14 20 21 
14 1 4 5 6 22 29 7 23 25 41 7 8 9 10 
14 1 4 5 6 22 29 7 23 25 41 7 15 9 17 
12 1 4 5 6 22 29 7 23 25 41 27 28 
8 1 4 5 6 34 35 27 28 
15 1 4 5 6 22 29 7 23 25 44 45 7 8 9 10 
13 1 4 5 6 22 29 7 23 25 44 45 27 28 
15 1 4 5 6 22 29 7 23 25 18 19 7 8 9 10 
15 1 4 5 6 22 29 7 23 25 18 19 7 15 9 17 
13 1 4 5 6 22 29 7 23 25 18 19 27 28 
16 1 4 5 6 22 29 7 23 25 18 19 29 7 20 9 21 
15 1 4 5 6 22 29 7 23 25 30 31 7 8 9 10 
15 1 4 5 6 22 29 7 23 25 30 31 7 15 9 17 
13 1 4 5 6 22 29 7 23 25 30 31 27 28 
16 1 4 5 6 22 29 7 23 25 30 31 29 7 20 9 21 
10 1 4 5 6 42 43 7 15 9 17 
8 1 4 5 6 34 35 20 21 
15 1 4 5 6 22 29 7 23 25 46 47 7 8 9 10 
13 1 4 5 6 22 29 7 23 25 46 47 27 28 
16 1 4 5 6 22 29 7 23 25 46 47 29 7 20 9 21 
18 1 4 5 6 22 29 7 23 25 22 29 7 23 25 7 8 9 10 
18 1 4 5 6 22 29 7 23 25 22 29 7 23 25 7 15 9 17 
16 1 4 5 6 22 29 7 23 25 22 29 7 23 25 27 28 
15 1 4 5 6 22 29 7 23 25 27 28 7 8 9 10 
15 1 4 5 6 22 29 7 23 25 27 28 7 15 9 17 
13 1 4 5 6 22 29 7 23 25 27 28 27 28 
15 1 4 5 6 22 29 7 23 25 13 32 7 8 9 10 
10 1 4 5 6 36 37 7 8 9 10 
15 1 4 5 6 22 29 7 23 25 13 32 7 15 9 17 
13 1 4 5 6 22 29 7 23 25 13 32 27 28 
14 1 4 5 6 22 29 7 23 25 33 7 8 9 10 
12 1 4 5 6 22 29 7 23 25 33 27 28 
15 1 4 5 6 22 29 7 23 25 34 35 7 8 9 10 
14 1 4 5 6 22 29 7 23 25 34 35 15 16 17 
13 1 4 5 6 22 29 7 23 25 34 35 27 28 
13 1 4 5 6 22 29 7 23 25 34 35 20 21 
15 1 4 5 6 22 29 7 23 25 36 37 7 8 9 10 
14 1 4 5 6 22 29 7 23 25 36 37 15 16 17 
9 1 4 5 6 36 37 15 16 17 
13 1 4 5 6 22 29 7 23 25 36 37 27 28 
16 1 4 5 6 22 29 7 23 25 36 37 29 7 20 9 21 
15 1 4 5 6 22 29 7 23 25 38 39 7 8 9 10 
15 1 4 5 6 22 29 7 23 25 38 39 7 15 9 17 
13 1 4 5 6 22 29 7 23 25 38 39 27 28 
14 1 4 5 6 22 29 7 23 25 40 7 8 9 10 
12 1 4 5 6 22 29 7 23 25 40 27 28 
12 1 4 5 6 27 28 30 31 7 8 9 10 
12 1 4 5 6 27 28 30 31 7 15 9 17 
10 1 4 5 6 27 28 30 31 27 28 
8 1 4 5 6 36 37 27 28 
13 1 4 5 6 27 28 30 31 29 7 20 9 21 
12 1 4 5 6 27 28 27 28 7 8 9 10 
12 1 4 5 6 27 28 27 28 7 15 9 17 
10 1 4 5 6 27 28 27 28 27 28 
12 1 4 5 6 27 28 38 39 7 8 9 10 
12 1 4 5 6 27 28 38 39 7 15 9 17 
10 1 4 5 6 27 28 38 39 27 28 
12 1 4 5 6 13 32 42 43 7 8 9 10 
10 1 4 5 6 13 32 42 43 27 28 
11 1 4 5 6 13 32 41 7 8 9 10 
11 1 4 5 6 36 37 29 7 20 9 21 
11 1 4 5 6 13 32 41 7 15 9 17 
9 1 4 5 6 13 32 41 27 28 
12 1 4 5 6 13 32 44 45 7 8 9 10 
10 1 4 5 6 13 32 44 45 27 28 
12 1 4 5 6 13 32 30 31 7 8 9 10 
12 1 4 5 6 13 32 30 31 7 15 9 17 
10 1 4 5 6 13 32 30 31 27 28 
13 1 4 5 6 13 32 30 31 29 7 20 9 21 
12 1 4 5 6 13 32 46 47 7 8 9 10 
10 1 4 5 6 13 32 46 47 27 28 
10 1 4 5 6 38 39 7 8 9 10 
13 1 4 5 6 13 32 46 47 29 7 20 9 21 
12 1 4 5 6 13 32 27 28 7 8 9 10 
12 1 4 5 6 13 32 27 28 7 15 9 17 
10 1 4 5 6 13 32 27 28 27 28 
12 1 4 5 6 13 32 13 32 7 8 9 10 
12 1 4 5 6 13 32 13 32 7 15 9 17 
10 1 4 5 6 13 32 13 32 27 28 
11 1 4 5 6 13 32 33 7 8 9 10 
9 1 4 5 6 13 32 33 27 28 
12 1 4 5 6 13 32 36 37 7 8 9 10 
10 1 4 5 6 38 39 7 15 9 17 
11 1 4 5 6 13 32 36 37 15 16 17 
10 1 4 5 6 13 32 36 37 27 28 
13 1 4 5 6 13 32 36 37 29 7 20 9 21 
12 1 4 5 6 13 32 38 39 7 8 9 10 
12 1 4 5 6 13 32 38 39 7 15 9 17 
10 1 4 5 6 13 32 38 39 27 28 
11 1 4 5 6 13 32 40 7 8 9 10 
9 1 4 5 6 13 32 40 27 28 
11 1 4 5 6 33 42 43 7 8 9 10 
9 1 4 5 6 33 42 43 27 28 
8 1 4 5 6 38 39 27 28 
11 1 4 5 6 33 44 45 7 8 9 10 
9 1 4 5 6 33 44 45 27 28 
11 1 4 5 6 33 46 47 7 8 9 10 
9 1 4 5 6 33 46 47 27 28 
12 1 4 5 6 33 46 47 29 7 20 9 21 
11 1 4 5 6 33 27 28 7 8 9 10 
11 1 4 5 6 33 27 28 7 15 9 17 
9 1 4 5 6 33 27 28 27 28 
10 1 4 5 6 33 33 7 8 9 10 
8 1 4 5 6 33 33 27 28 
11 1 4 5 6 38 39 29 7 20 9 21 
10 1 4 5 6 33 40 7 8 9 10 
8 1 4 5 6 33 40 27 28 
12 1 4 5 6 34 35 42 43 7 8 9 10 
10 1 4 5 6 34 35 42 43 27 28 
14 1 4 5 6 34 35 11 12 13 14 7 8 9 10 
13 1 4 5 6 34 35 11 12 13 14 15 16 17 
12 1 4 5 6 34 35 11 12 13 14 27 28 
12 1 4 5 6 34 35 11 12 13 14 20 21 
11 1 4 5 6 34 35 41 7 8 9 10 
10 1 4 5 6 34 35 41 15 16 17 
9 1 4 5 6 40 7 8 9 10 
9 1 4 5 6 34 35 41 27 28 
12 1 4 5 6 34 35 44 45 7 8 9 10 
10 1 4 5 6 34 35 44 45 27 28 
12 1 4 5 6 34 35 18 19 7 8 9 10 
11 1 4 5 6 34 35 18 19 15 16 17 
10 1 4 5 6 34 35 18 19 27 28 
10 1 4 5 6 34 35 18 19 20 21 
12 1 4 5 6 34 35 30 31 7 8 9 10 
11 1 4 5 6 34 35 30 31 15 16 17 
10 1 4 5 6 34 35 30 31 27 28 
8 1 4 5 6 42 43 27 28 
9 1 4 5 6 40 7 15 9 17 
10 1 4 5 6 34 35 30 31 20 21 
12 1 4 5 6 34 35 46 47 7 8 9 10 
10 1 4 5 6 34 35 46 47 27 28 
10 1 4 5 6 34 35 46 47 20 21 
15 1 4 5 6 34 35 22 23 26 24 25 7 8 9 10 
14 1 4 5 6 34 35 22 23 24 25 7 8 9 10 
14 1 4 5 6 34 35 22 23 26 24 25 15 16 17 
13 1 4 5 6 34 35 22 23 24 25 15 16 17 
13 1 4 5 6 34 35 22 23 26 24 25 27 28 
12 1 4 5 6 34 35 22 23 24 25 27 28 
7 1 4 5 6 40 27 28 
11 1 4 5 6 34 35 15 16 17 8 10 
12 1 4 5 6 34 35 15 16 17 15 16 17 
13 1 4 5 6 34 35 15 16 17 7 27 9 28 
14 1 4 5 6 34 35 15 16 17 29 7 20 9 21 
12 1 4 5 6 34 35 27 28 7 8 9 10 
11 1 4 5 6 34 35 27 28 15 16 17 
10 1 4 5 6 34 35 27 28 27 28 
12 1 4 5 6 34 35 13 32 7 8 9 10 
11 1 4 5 6 34 35 13 32 15 16 17 
10 1 4 5 6 34 35 13 32 27 28 
10 1 4 5 6 40 29 7 20 9 21 
11 1 4 5 6 34 35 33 7 8 9 10 
9 1 4 5 6 34 35 33 27 28 
12 1 4 5 6 34 35 34 35 7 8 9 10 
11 1 4 5 6 34 35 34 35 15 16 17 
10 1 4 5 6 34 35 34 35 27 28 
10 1 4 5 6 34 35 34 35 20 21 
12 1 4 5 6 34 35 36 37 7 8 9 10 
11 1 4 5 6 34 35 36 37 15 16 17 
10 1 4 5 6 34 35 36 37 27 28 
10 1 4 5 6 34 35 36 37 20 21 
9 1 4 5 6 29 7 20 9 21 
12 1 4 5 6 34 35 38 39 7 8 9 10 
11 1 4 5 6 34 35 38 39 15 16 17 
10 1 4 5 6 34 35 38 39 27 28 
11 1 4 5 6 34 35 40 7 8 9 10 
9 1 4 5 6 34 35 40 27 28 
12 1 4 5 6 34 35 20 21 7 8 9 10 
11 1 4 5 6 34 35 20 21 15 16 17 
10 1 4 5 6 34 35 20 21 27 28 
10 1 4 5 6 34 35 20 21 20 21 
12 1 4 5 6 38 39 42 43 7 8 9 10 
9 1 4 5 6 29 7 20 9 21 
10 1 4 5 6 38 39 42 43 27 28 
12 1 4 5 6 38 39 44 45 7 8 9 10 
10 1 4 5 6 38 39 44 45 27 28 
12 1 4 5 6 38 39 30 31 7 8 9 10 
12 1 4 5 6 38 39 30 31 7 15 9 17 
10 1 4 5 6 38 39 30 31 27 28 
13 1 4 5 6 38 39 30 31 29 7 20 9 21 
12 1 4 5 6 38 39 46 47 7 8 9 10 
10 1 4 5 6 38 39 46 47 27 28 
13 1 4 5 6 38 39 46 47 29 7 20 9 21 
9 1 4 5 6 29 7 20 9 21 
15 1 4 5 6 38 39 22 29 7 23 25 7 8 9 10 
15 1 4 5 6 38 39 22 29 7 23 25 7 15 9 17 
13 1 4 5 6 38 39 22 29 7 23 25 27 28 
12 1 4 5 6 38 39 27 28 7 8 9 10 
12 1 4 5 6 38 39 27 28 7 15 9 17 
10 1 4 5 6 38 39 27 28 27 28 
11 1 4 5 6 38 39 33 7 8 9 10 
9 1 4 5 6 38 39 33 27 28 
12 1 4 5 6 38 39 38 39 7 8 9 10 
12 1 4 5 6 38 39 38 39 7 15 9 17 
9 1 4 5 6 29 7 20 9 21 
10 1 4 5 6 38 39 38 39 27 28 
11 1 4 5 6 38 39 40 7 8 9 10 
9 1 4 5 6 38 39 40 27 28 
11 1 4 5 6 40 42 43 7 8 9 10 
9 1 4 5 6 40 42 43 27 28 
11 1 4 5 6 40 44 45 7 8 9 10 
9 1 4 5 6 40 44 45 27 28 
11 1 4 5 6 40 27 28 7 8 9 10 
11 1 4 5 6 40 27 28 7 15 9 17 
9 1 4 5 6 40 27 28 27 28 
14 1 4 5 6 11 12 13 14 42 43 7 8 9 10 
10 1 4 5 6 40 40 7 8 9 10 
8 1 4 5 6 40 40 27 28 
14 1 4 5 6 42 43 42 43 42 43 7 8 9 10 
12 1 4 5 6 42 43 42 43 42 43 27 28 
16 1 4 5 6 42 43 42 43 11 12 13 14 7 8 9 10 
15 1 4 5 6 42 43 42 43 11 12 13 14 15 16 17 
14 1 4 5 6 42 43 42 43 11 12 13 14 27 28 
14 1 4 5 6 42 43 42 43 11 12 13 14 20 21 
17 1 4 5 6 42 43 42 43 22 29 7 23 25 7 8 9 10 
17 1 4 5 6 42 43 42 43 22 29 7 23 25 7 15 9 17 
13 1 4 5 6 11 12 13 14 42 43 15 16 17 
15 1 4 5 6 42 43 42 43 22 29 7 23 25 27 28 
14 1 4 5 6 42 43 42 43 27 28 7 8 9 10 
14 1 4 5 6 42 43 42 43 27 28 7 15 9 17 
12 1 4 5 6 42 43 42 43 27 28 27 28 
14 1 4 5 6 42 43 42 43 34 35 7 8 9 10 
13 1 4 5 6 42 43 42 43 34 35 15 16 17 
12 1 4 5 6 42 43 42 43 34 35 27 28 
12 1 4 5 6 42 43 42 43 34 35 20 21 
16 1 4 5 6 42 43 11 12 13 14 42 43 7 8 9 10 
14 1 4 5 6 42 43 11 12 13 14 42 43 27 28 
12 1 4 5 6 11 12 13 14 42 43 27 28 
18 1 4 5 6 42 43 11 12 13 14 11 12 13 14 7 8 9 10 
17 1 4 5 6 42 43 11 12 13 14 11 12 13 14 15 16 17 
16 1 4 5 6 42 43 11 12 13 14 11 12 13 14 27 28 
16 1 4 5 6 42 43 11 12 13 14 11 12 13 14 20 21 
15 1 4 5 6 42 43 11 12 13 14 41 7 8 9 10 
14 1 4 5 6 42 43 11 12 13 14 41 15 16 17 
13 1 4 5 6 42 43 11 12 13 14 41 27 28 
16 1 4 5 6 42 43 11 12 13 14 44 45 7 8 9 10 
14 1 4 5 6 42 43 11 12 13 14 44 45 27 28 
16 1 4 5 6 42 43 11 12 13 14 18 19 7 8 9 10 
11 1 4 5 6 42 43 29 7 20 9 21 
12 1 4 5 6 11 12 13 14 42 43 20 21 
15 1 4 5 6 42 43 11 12 13 14 18 19 15 16 17 
14 1 4 5 6 42 43 11 12 13 14 18 19 27 28 
14 1 4 5 6 42 43 11 12 13 14 18 19 20 21 
16 1 4 5 6 42 43 11 12 13 14 30 31 7 8 9 10 
15 1 4 5 6 42 43 11 12 13 14 30 31 15 16 17 
14 1 4 5 6 42 43 11 12 13 14 30 31 27 28 
14 1 4 5 6 42 43 11 12 13 14 30 31 20 21 
16 1 4 5 6 42 43 11 12 13 14 46 47 7 8 9 10 
14 1 4 5 6 42 43 11 12 13 14 46 47 27 28 
14 1 4 5 6 42 43 11 12 13 14 46 47 20 21 
16 1 4 5 6 11 12 13 14 11 12 13 14 7 8 9 10 
19 1 4 5 6 42 43 11 12 13 14 22 23 26 24 25 7 8 9 10 
18 1 4 5 6 42 43 11 12 13 14 22 23 24 25 7 8 9 10 
18 1 4 5 6 42 43 11 12 13 14 22 23 26 24 25 15 16 17 
17 1 4 5 6 42 43 11 12 13 14 22 23 24 25 15 16 17 
17 1 4 5 6 42 43 11 12 13 14 22 23 26 24 25 27 28 
16 1 4 5 6 42 43 11 12 13 14 22 23 24 25 27 28 
15 1 4 5 6 42 43 11 12 13 14 15 16 17 8 10 
16 1 4 5 6 42 43 11 12 13 14 15 16 17 15 16 17 
17 1 4 5 6 42 43 11 12 13 14 15 16 17 7 27 9 28 
18 1 4 5 6 42 43 11 12 13 14 15 16 17 29 7 20 9 21 
15 1 4 5 6 11 12 13 14 11 12 13 14 15 16 17 
16 1 4 5 6 42 43 11 12 13 14 27 28 7 8 9 10 
15 1 4 5 6 42 43 11 12 13 14 27 28 15 16 17 
14 1 4 5 6 42 43 11 12 13 14 27 28 27 28 
16 1 4 5 6 42 43 11 12 13 14 13 32 7 8 9 10 
15 1 4 5 6 42 43 11 12 13 14 13 32 15 16 17 
14 1 4 5 6 42 43 11 12 13 14 13 32 27 28 
15 1 4 5 6 42 43 11 12 13 14 33 7 8 9 10 
13 1 4 5 6 42 43 11 12 13 14 33 27 28 
16 1 4 5 6 42 43 11 12 13 14 34 35 7 8 9 10 
15 1 4 5 6 42 43 11 12 13 14 34 35 15 16 17 
14 1 4 5 6 11 12 13 14 11 12 13 14 27 28 
14 1 4 5 6 42 43 11 12 13 14 34 35 27 28 
14 1 4 5 6 42 43 11 12 13 14 34 35 20 21 
16 1 4 5 6 42 43 11 12 13 14 36 37 7 8 9 10 
15 1 4 5 6 42 43 11 12 13 14 36 37 15 16 17 
14 1 4 5 6 42 43 11 12 13 14 36 37 27 28 
14 1 4 5 6 42 43 11 12 13 14 36 37 20 21 
16 1 4 5 6 42 43 11 12 13 14 38 39 7 8 9 10 
15 1 4 5 6 42 43 11 12 13 14 38 39 15 16 17 
14 1 4 5 6 42 43 11 12 13 14 38 39 27 28 
15 1 4 5 6 42 43 11 12 13 14 40 7 8 9 10 
14 1 4 5 6 11 12 13 14 11 12 13 14 20 21 
13 1 4 5 6 42 43 11 12 13 14 40 27 28 
16 1 4 5 6 42 43 11 12 13 14 20 21 7 8 9 10 
15 1 4 5 6 42 43 11 12 13 14 20 21 15 16 17 
14 1 4 5 6 42 43 11 12 13 14 20 21 27 28 
14 1 4 5 6 42 43 11 12 13 14 20 21 20 21 
17 1 4 5 6 42 43 22 29 7 23 25 42 43 7 8 9 10 
15 1 4 5 6 42 43 22 29 7 23 25 42 43 27 28 
19 1 4 5 6 42 43 22 29 7 23 25 11 12 13 14 7 8 9 10 
18 1 4 5 6 42 43 22 29 7 23 25 11 12 13 14 15 16 17 
17 1 4 5 6 42 43 22 29 7 23 25 11 12 13 14 27 28 
12 1 4 5 6 11 12 13 14 7 8 9 10 
17 1 4 5 6 42 43 22 29 7 23 25 11 12 13 14 20 21 
16 1 4 5 6 42 43 22 29 7 23 25 41 7 8 9 10 
16 1 4 5 6 42 43 22 29 7 23 25 41 7 15 9 17 
14 1 4 5 6 42 43 22 29 7 23 25 41 27 28 
17 1 4 5 6 42 43 22 29 7 23 25 44 45 7 8 9 10 
15 1 4 5 6 42 43 22 29 7 23 25 44 45 27 28 
17 1 4 5 6 42 43 22 29 7 23 25 18 19 7 8 9 10 
17 1 4 5 6 42 43 22 29 7 23 25 18 19 7 15 9 17 
15 1 4 5 6 42 43 22 29 7 23 25 18 19 27 28 
18 1 4 5 6 42 43 22 29 7 23 25 18 19 29 7 20 9 21 
12 1 4 5 6 11 12 13 14 7 8 9 10 
17 1 4 5 6 42 43 22 29 7 23 25 30 31 7 8 9 10 
17 1 4 5 6 42 43 22 29 7 23 25 30 31 7 15 9 17 
15 1 4 5 6 42 43 22 29 7 23 25 30 31 27 28 
18 1 4 5 6 42 43 22 29 7 23 25 30 31 29 7 20 9 21 
17 1 4 5 6 42 43 22 29 7 23 25 46 47 7 8 9 10 
15 1 4 5 6 42 43 22 29 7 23 25 46 47 27 28 
18 1 4 5 6 42 43 22 29 7 23 25 46 47 29 7 20 9 21 
20 1 4 5 6 42 43 22 29 7 23 25 22 29 7 23 25 7 8 9 10 
20 1 4 5 6 42 43 22 29 7 23 25 22 29 7 23 25 7 15 9 17 
18 1 4 5 6 42 43 22 29 7 23 25 22 29 7 23 25 27 28 
12 1 4 5 6 11 12 13 14 7 8 9 10 
17 1 4 5 6 42 43 22 29 7 23 25 27 28 7 8 9 10 
17 1 4 5 6 42 43 22 29 7 23 25 27 28 7 15 9 17 
15 1 4 5 6 42 43 22 29 7 23 25 27 28 27 28 
17 1 4 5 6 42 43 22 29 7 23 25 13 32 7 8 9 10 
17 1 4 5 6 42 43 22 29 7 23 25 13 32 7 15 9 17 
15 1 4 5 6 42 43 22 29 7 23 25 13 32 27 28 
16 1 4 5 6 42 43 22 29 7 23 25 33 7 8 9 10 
14 1 4 5 6 42 43 22 29 7 23 25 33 27 28 
17 1 4 5 6 42 43 22 29 7 23 25 34 35 7 8 9 10 
16 1 4 5 6 42 43 22 29 7 23 25 34 35 15 16 17 
12 1 4 5 6 11 12 13 14 7 8 9 10 
15 1 4 5 6 42 43 22 29 7 23 25 34 35 27 28 
15 1 4 5 6 42 43 22 29 7 23 25 34 35 20 21 
17 1 4 5 6 42 43 22 29 7 23 25 36 37 7 8 9 10 
16 1 4 5 6 42 43 22 29 7 23 25 36 37 15 16 17 
15 1 4 5 6 42 43 22 29 7 23 25 36 37 27 28 
18 1 4 5 6 42 43 22 29 7 23 25 36 37 29 7 20 9 21 
17 1 4 5 6 42 43 22 29 7 23 25 38 39 7 8 9 10 
17 1 4 5 6 42 43 22 29 7 23 25 38 39 7 15 9 17 
15 1 4 5 6 42 43 22 29 7 23 25 38 39 27 28 
16 1 4 5 6 42 43 22 29 7 23 25 40 7 8 9 10 
13 1 4 5 6 11 12 13 14 41 7 8 9 10 
14 1 4 5 6 42 43 22 29 7 23 25 40 27 28 
14 1 4 5 6 42 43 27 28 30 31 7 8 9 10 
14 1 4 5 6 42 43 27 28 30 31 7 15 9 17 
12 1 4 5 6 42 43 27 28 30 31 27 28 
15 1 4 5 6 42 43 27 28 30 31 29 7 20 9 21 
14 1 4 5 6 42 43 27 28 27 28 7 8 9 10 
14 1 4 5 6 42 43 27 28 27 28 7 15 9 17 
12 1 4 5 6 42 43 27 28 27 28 27 28 
14 1 4 5 6 42 43 27 28 38 39 7 8 9 10 
14 1 4 5 6 42 43 27 28 38 39 7 15 9 17 
12 1 4 5 6 11 12 13 14 7 8 9 10 
12 1 4 5 6 11 12 13 14 41 15 16 17 
12 1 4 5 6 42 43 27 28 38 39 27 28 
14 1 4 5 6 42 43 34 35 42 43 7 8 9 10 
12 1 4 5 6 42 43 34 35 42 43 27 28 
16 1 4 5 6 42 43 34 35 11 12 13 14 7 8 9 10 
15 1 4 5 6 42 43 34 35 11 12 13 14 15 16 17 
14 1 4 5 6 42 43 34 35 11 12 13 14 27 28 
14 1 4 5 6 42 43 34 35 11 12 13 14 20 21 
13 1 4 5 6 42 43 34 35 41 7 8 9 10 
12 1 4 5 6 42 43 34 35 41 15 16 17 
11 1 4 5 6 42 43 34 35 41 27 28 
11 1 4 5 6 11 12 13 14 41 27 28 
14 1 4 5 6 42 43 34 35 44 45 7 8 9 10 
12 1 4 5 6 42 43 34 35 44 45 27 28 
14 1 4 5 6 42 43 34 35 18 19 7 8 9 10 
13 1 4 5 6 42 43 34 35 18 19 15 16 17 
12 1 4 5 6 42 43 34 35 18 19 27 28 
12 1 4 5 6 42 43 34 35 18 19 20 21 
14 1 4 5 6 42 43 34 35 30 31 7 8 9 10 
13 1 4 5 6 42 43 34 35 30 31 15 16 17 
12 1 4 5 6 42 43 34 35 30 31 27 28 
12 1 4 5 6 42 43 34 35 30 31 20 21 
11 1 4 5 6 11 12 13 14 41 20 21 
14 1 4 5 6 42 43 34 35 46 47 7 8 9 10 
12 1 4 5 6 42 43 34 35 46 47 27 28 
12 1 4 5 6 42 43 34 35 46 47 20 21 
17 1 4 5 6 42 43 34 35 22 23 26 24 25 7 8 9 10 
16 1 4 5 6 42 43 34 35 22 23 24 25 7 8 9 10 
16 1 4 5 6 42 43 34 35 22 23 26 24 25 15 16 17 
15 1 4 5 6 42 43 34 35 22 23 24 25 15 16 17 
15 1 4 5 6 42 43 34 35 22 23 26 24 25 27 28 
14 1 4 5 6 42 43 34 35 22 23 24 25 27 28 
13 1 4 5 6 42 43 34 35 15 16 17 8 10 
14 1 4 5 6 11 12 13 14 44 45 7 8 9 10 
14 1 4 5 6 42 43 34 35 15 16 17 15 16 17 
15 1 4 5 6 42 43 34 35 15 16 17 7 27 9 28 
16 1 4 5 6 42 43 34 35 15 16 17 29 7 20 9 21 
14 1 4 5 6 42 43 34 35 27 28 7 8 9 10 
13 1 4 5 6 42 43 34 35 27 28 15 16 17 
12 1 4 5 6 42 43 34 35 27 28 27 28 
14 1 4 5 6 42 43 34 35 13 32 7 8 9 10 
13 1 4 5 6 42 43 34 35 13 32 15 16 17 
12 1 4 5 6 42 43 34 35 13 32 27 28 
13 1 4 5 6 42 43 34 35 33 7 8 9 10 
13 1 4 5 6 11 12 13 14 44 45 15 16 17 
11 1 4 5 6 42 43 34 35 33 27 28 
14 1 4 5 6 42 43 34 35 34 35 7 8 9 10 
13 1 4 5 6 42 43 34 35 34 35 15 16 17 
12 1 4 5 6 42 43 34 35 34 35 27 28 
12 1 4 5 6 42 43 34 35 34 35 20 21 
14 1 4 5 6 42 43 34 35 36 37 7 8 9 10 
13 1 4 5 6 42 43 34 35 36 37 15 16 17 
12 1 4 5 6 42 43 34 35 36 37 27 28 
12 1 4 5 6 42 43 34 35 36 37 20 21 
14 1 4 5 6 42 43 34 35 38 39 7 8 9 10 
12 1 4 5 6 11 12 13 14 44 45 27 28 
13 1 4 5 6 42 43 34 35 38 39 15 16 17 
12 1 4 5 6 42 43 34 35 38 39 27 28 
13 1 4 5 6 42 43 34 35 40 7 8 9 10 
11 1 4 5 6 42 43 34 35 40 27 28 
14 1 4 5 6 42 43 34 35 20 21 7 8 9 10 
13 1 4 5 6 42 43 34 35 20 21 15 16 17 
12 1 4 5 6 42 43 34 35 20 21 27 28 
12 1 4 5 6 42 43 34 35 20 21 20 21 
16 1 4 5 6 11 12 13 14 42 43 42 43 7 8 9 10 
14 1 4 5 6 11 12 13 14 42 43 42 43 27 28 
12 1 4 5 6 11 12 13 14 44 45 20 21 
18 1 4 5 6 11 12 13 14 42 43 11 12 13 14 7 8 9 10 
17 1 4 5 6 11 12 13 14 42 43 11 12 13 14 15 16 17 
16 1 4 5 6 11 12 13 14 42 43 11 12 13 14 27 28 
16 1 4 5 6 11 12 13 14 42 43 11 12 13 14 20 21 
19 1 4 5 6 11 12 13 14 42 43 22 23 26 24 25 7 8 9 10 
18 1 4 5 6 11 12 13 14 42 43 22 23 24 25 7 8 9 10 
18 1 4 5 6 11 12 13 14 42 43 22 23 26 24 25 15 16 17 
17 1 4 5 6 11 12 13 14 42 43 22 23 24 25 15 16 17 
17 1 4 5 6 11 12 13 14 42 43 22 23 26 24 25 27 28 
16 1 4 5 6 11 12 13 14 42 43 22 23 24 25 27 28 
14 1 4 5 6 11 12 13 14 18 19 7 8 9 10 
16 1 4 5 6 11 12 13 14 42 43 27 28 7 8 9 10 
15 1 4 5 6 11 12 13 14 42 43 27 28 15 16 17 
14 1 4 5 6 11 12 13 14 42 43 27 28 27 28 
16 1 4 5 6 11 12 13 14 42 43 34 35 7 8 9 10 
15 1 4 5 6 11 12 13 14 42 43 34 35 15 16 17 
14 1 4 5 6 11 12 13 14 42 43 34 35 27 28 
14 1 4 5 6 11 12 13 14 42 43 34 35 20 21 
18 1 4 5 6 11 12 13 14 11 12 13 14 42 43 7 8 9 10 
16 1 4 5 6 11 12 13 14 11 12 13 14 42 43 27 28 
20 1 4 5 6 11 12 13 14 11 12 13 14 11 12 13 14 7 8 9 10 
13 1 4 5 6 11 12 13 14 18 19 15 16 17 
19 1 4 5 6 11 12 13 14 11 12 13 14 11 12 13 14 15 16 17 
18 1 4 5 6 11 12 13 14 11 12 13 14 11 12 13 14 27 28 
18 1 4 5 6 11 12 13 14 11 12 13 14 11 12 13 14 20 21 
17 1 4 5 6 11 12 13 14 11 12 13 14 41 7 8 9 10 
16 1 4 5 6 11 12 13 14 11 12 13 14 41 15 16 17 
15 1 4 5 6 11 12 13 14 11 12 13 14 41 27 28 
18 1 4 5 6 11 12 13 14 11 12 13 14 44 45 7 8 9 10 
16 1 4 5 6 11 12 13 14 11 12 13 14 44 45 27 28 
18 1 4 5 6 11 12 13 14 11 12 13 14 18 19 7 8 9 10 
17 1 4 5 6 11 12 13 14 11 12 13 14 18 19 15 16 17 
12 1 4 5 6 11 12 13 14 18 19 27 28 
16 1 4 5 6 11 12 13 14 11 12 13 14 18 19 27 28 
16 1 4 5 6 11 12 13 14 11 12 13 14 18 19 20 21 
18 1 4 5 6 11 12 13 14 11 12 13 14 30 31 7 8 9 10 
17 1 4 5 6 11 12 13 14 11 12 13 14 30 31 15 16 17 
16 1 4 5 6 11 12 13 14 11 12 13 14 30 31 27 28 
16 1 4 5 6 11 12 13 14 11 12 13 14 30 31 20 21 
18 1 4 5 6 11 12 13 14 11 12 13 14 46 47 7 8 9 10 
16 1 4 5 6 11 12 13 14 11 12 13 14 46 47 27 28 
16 1 4 5 6 11 12 13 14 11 12 13 14 46 47 20 21 
21 1 4 5 6 11 12 13 14 11 12 13 14 22 23 26 24 25 7 8 9 10 
