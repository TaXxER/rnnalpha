1050 17
22 1 2 3 4 5 6 7 8 9 3 2 2 3 2 3 3 2 2 3 3 2 10 
12 1 5 3 4 2 6 7 8 9 3 3 10 
14 1 5 6 2 3 7 8 9 9 2 3 2 3 10 
13 1 5 6 3 4 2 7 8 9 2 3 10 11 
8 1 5 6 7 3 2 4 8 
10 1 5 6 2 3 4 8 7 9 10 
12 1 5 6 7 8 4 3 2 9 2 3 10 
13 1 5 6 3 4 2 12 9 3 2 3 9 13 
11 1 5 6 8 2 3 4 9 2 3 10 
11 1 5 6 3 2 4 7 8 9 3 10 
16 1 5 6 4 3 2 8 9 2 3 9 7 3 2 10 11 
15 1 5 6 2 3 4 7 8 9 2 2 2 3 10 11 
3 1 5 6 
12 1 5 6 3 4 2 9 7 8 3 2 10 
11 1 5 6 7 3 2 4 8 9 10 11 
3 1 5 6 
3 1 5 6 
5 1 5 6 3 2 
19 1 5 6 2 3 4 7 8 9 12 4 2 3 9 2 3 2 10 11 
10 1 5 6 7 8 3 4 2 9 13 
11 1 5 6 2 9 2 2 2 2 3 13 
21 1 5 6 7 2 4 3 8 12 4 3 2 4 4 3 2 9 2 3 10 11 
11 1 5 6 7 4 2 3 8 9 3 10 
13 1 5 2 3 4 6 2 3 4 9 3 10 11 
8 1 5 6 8 3 4 2 7 
10 1 5 6 2 4 3 12 9 9 10 
8 1 5 6 2 4 3 7 8 
13 1 5 6 7 8 4 3 2 9 3 2 10 11 
8 1 5 6 7 8 3 4 2 
12 1 5 6 3 2 4 8 9 7 2 3 14 
15 1 5 6 2 3 4 7 8 9 9 2 3 3 10 11 
8 1 5 3 4 2 6 7 8 
12 1 5 6 7 8 3 2 4 9 3 2 10 
11 1 5 2 3 4 6 9 9 2 3 10 
8 7 1 5 6 4 3 2 8 
14 1 6 8 5 2 4 3 9 9 3 4 2 10 11 
16 1 5 6 7 8 3 4 2 9 2 3 2 3 3 2 10 
5 1 5 6 2 3 
14 1 5 6 4 2 3 7 8 9 2 3 3 2 10 
24 1 5 6 8 7 2 3 4 9 9 2 3 3 2 2 2 2 2 3 4 2 3 2 14 
11 1 5 6 7 8 4 3 2 2 3 4 
6 1 5 6 2 3 4 
14 1 5 6 7 2 4 3 8 9 3 2 3 2 15 
3 1 5 6 
14 1 5 6 7 3 4 2 8 9 3 2 3 10 11 
10 1 5 6 3 2 9 3 2 3 10 
11 1 5 6 4 2 3 7 8 9 4 10 
13 1 5 6 3 4 2 7 8 9 3 2 9 10 
8 1 5 6 3 9 9 10 11 
3 1 5 6 
6 1 5 6 2 3 4 
8 1 5 6 3 4 2 7 8 
8 1 5 6 3 4 2 7 8 
6 1 5 6 3 4 2 
14 1 5 6 3 4 2 7 8 9 9 3 2 3 10 
12 1 5 6 3 4 2 7 8 9 2 3 10 
8 1 5 6 2 3 4 7 8 
8 1 5 6 7 8 3 2 4 
13 1 2 4 3 5 6 7 8 9 2 3 10 11 
15 1 5 6 3 4 2 7 8 9 3 2 9 2 3 10 
14 1 2 3 4 5 6 7 8 9 2 9 3 2 10 
8 1 5 6 3 4 2 7 8 
11 1 5 6 4 3 2 8 7 9 10 11 
19 1 5 4 3 2 6 7 8 9 9 3 2 2 3 3 2 2 3 13 
3 1 5 6 
21 1 5 6 2 4 3 7 8 9 3 2 4 9 3 2 3 3 2 3 2 10 
16 1 5 3 4 2 6 7 8 9 3 2 2 3 2 3 10 
16 1 5 6 7 3 4 2 8 9 2 3 2 3 2 10 11 
16 1 5 6 7 3 4 2 8 9 3 2 2 3 2 10 11 
7 1 5 6 2 3 9 10 
14 1 5 6 7 8 2 3 4 9 3 9 3 10 11 
9 1 5 6 2 4 3 9 10 11 
9 1 5 6 7 3 4 2 8 9 
13 1 5 6 2 3 4 8 9 9 3 2 10 11 
5 1 5 6 3 2 
11 1 5 6 2 4 3 7 8 9 4 13 
15 1 5 6 3 4 2 8 7 9 9 3 2 2 3 10 
16 1 5 6 2 4 3 8 9 7 2 3 2 3 2 10 11 
13 1 5 6 2 4 3 7 8 9 3 2 10 11 
5 1 5 6 2 3 
14 1 5 6 7 8 3 2 4 9 9 3 2 15 11 
12 1 5 6 4 2 3 7 8 9 3 10 11 
17 1 5 6 4 2 3 7 8 9 3 2 2 3 2 3 2 10 
7 1 5 6 2 3 9 10 
12 1 5 6 7 8 2 3 4 9 3 2 10 
5 1 5 6 2 3 
12 5 1 6 7 8 2 3 4 9 2 10 11 
15 1 5 6 7 8 2 3 4 9 3 2 3 2 10 11 
13 1 5 6 2 4 3 7 8 9 3 2 3 10 
21 1 5 6 3 4 2 8 9 9 3 3 2 3 3 2 3 2 3 2 10 11 
14 1 5 6 7 2 3 4 8 9 2 3 2 10 11 
7 1 5 6 2 3 8 7 
22 1 5 6 7 8 2 3 3 2 4 12 3 4 2 2 3 4 9 2 3 10 11 
5 1 5 6 2 3 
15 1 5 6 2 3 4 7 8 9 3 2 3 2 3 10 
13 1 5 6 3 2 7 8 9 9 3 3 10 11 
9 1 5 6 3 4 2 8 7 4 
24 1 7 5 6 8 3 4 2 12 3 4 2 3 2 4 4 3 2 2 3 4 9 10 11 
32 1 5 6 7 2 3 8 9 12 4 3 2 2 3 4 4 2 4 3 2 4 4 2 4 3 9 2 3 2 3 10 11 
13 1 5 6 4 2 3 8 7 9 3 2 3 10 
12 7 1 5 6 4 3 2 8 9 9 10 11 
8 1 5 6 7 8 4 2 3 
9 3 2 1 5 2 3 6 7 8 
10 1 4 3 2 5 6 4 4 7 8 
29 1 5 6 4 3 2 7 8 9 12 2 4 3 4 2 3 2 3 4 3 4 2 9 3 2 2 3 10 11 
12 1 5 7 6 3 4 2 8 9 2 3 10 
8 1 5 6 2 4 3 7 8 
8 1 5 6 2 3 4 9 13 
33 1 5 6 2 3 4 7 8 9 2 9 2 2 3 3 3 2 2 2 2 2 3 9 9 2 2 3 3 2 3 2 10 11 
11 1 5 6 3 2 4 7 8 3 2 4 
14 1 5 6 2 4 3 7 8 9 2 3 2 3 14 
32 1 5 2 3 4 6 7 8 12 12 2 3 4 2 3 4 2 2 3 4 4 3 4 2 4 2 3 2 4 3 9 10 
3 1 5 6 
14 1 4 2 3 5 6 7 8 9 9 2 3 10 11 
17 6 1 5 2 3 4 7 8 12 4 3 3 4 2 9 10 11 
14 1 5 6 7 3 4 2 8 9 2 3 2 3 10 
15 1 5 3 4 2 6 7 8 9 2 3 3 2 10 11 
16 1 5 6 3 2 4 8 9 9 7 3 2 2 3 2 10 
118 1 3 2 5 6 7 8 12 4 3 2 4 4 2 3 3 2 4 2 3 4 3 4 2 2 3 4 2 4 3 3 4 2 2 3 4 3 2 4 3 2 4 4 2 3 4 3 2 2 3 4 4 2 3 3 2 4 2 3 4 3 4 2 4 3 2 2 3 4 4 3 2 4 2 3 2 3 4 2 4 3 3 2 4 3 4 2 2 3 2 4 2 3 4 2 4 3 4 2 3 3 4 2 2 3 4 4 4 3 2 2 2 3 4 3 4 2 13 
9 1 2 4 3 5 6 7 8 2 
12 1 5 6 3 4 2 8 9 9 3 2 13 
7 1 5 6 2 3 7 8 
14 1 5 3 4 2 6 8 7 9 2 3 2 3 10 
16 1 5 6 2 3 8 9 4 9 9 7 2 3 3 2 13 
31 1 5 6 3 4 2 7 8 9 4 2 3 9 2 3 3 2 2 3 3 2 3 3 3 2 3 2 3 3 15 11 
11 1 2 4 3 5 6 8 9 9 7 10 
3 1 5 6 
10 1 7 5 6 8 3 4 2 9 10 
8 1 5 6 4 2 3 7 8 
7 1 5 6 3 2 9 10 
18 1 5 6 2 3 4 7 8 9 2 3 12 2 4 3 9 10 11 
15 1 5 6 2 3 4 8 7 9 2 9 3 2 10 11 
11 1 5 6 2 4 3 7 8 9 9 10 
5 1 5 6 3 2 
7 1 5 6 2 3 9 10 
17 1 5 2 4 3 6 9 3 2 3 2 3 2 3 2 10 11 
15 1 5 6 2 4 3 7 8 9 9 2 3 3 2 10 
17 1 5 6 3 4 2 7 8 9 2 3 9 2 3 3 3 10 
7 1 5 6 2 3 9 10 
16 1 5 6 2 3 4 8 7 9 9 2 3 3 2 10 11 
16 1 5 6 3 4 2 8 7 9 2 3 9 2 3 10 11 
12 1 5 6 3 2 4 8 7 9 2 3 13 
15 1 5 3 4 2 6 7 8 9 3 2 3 2 10 11 
5 1 5 6 3 2 
3 1 5 6 
8 1 5 6 7 8 3 2 4 
21 1 5 6 2 4 3 7 8 12 3 4 2 9 3 2 3 2 2 3 10 11 
8 1 5 6 7 3 2 4 8 
10 1 5 6 7 3 4 2 8 9 10 
5 1 5 3 2 6 
19 1 5 6 7 8 2 3 4 9 3 2 9 3 2 2 3 2 3 10 
19 1 5 6 4 3 2 7 8 12 2 3 4 4 3 2 3 4 2 10 
17 1 5 3 4 2 6 12 4 2 3 4 2 3 4 9 10 11 
8 1 5 6 7 8 2 4 3 
13 1 5 6 4 2 3 7 8 9 9 2 3 10 
16 1 5 6 2 4 3 7 8 9 2 2 3 2 2 3 13 
17 1 3 2 5 6 4 7 8 9 3 2 2 3 3 2 10 11 
13 1 5 6 7 2 3 4 8 9 2 3 10 11 
27 1 5 6 4 3 2 8 9 3 2 3 2 2 3 2 3 3 2 2 3 2 3 3 3 2 10 11 
5 1 5 3 2 6 
14 1 4 3 2 5 6 8 7 9 2 3 2 3 10 
8 1 5 6 3 2 4 7 8 
59 1 5 6 2 3 4 7 8 12 2 3 4 3 4 2 4 2 3 2 3 4 2 3 4 2 4 3 2 4 2 3 2 3 4 9 2 3 3 2 3 2 2 2 2 3 3 2 3 2 2 3 3 2 3 2 2 3 10 11 
13 1 5 6 7 2 3 4 8 9 9 2 3 10 
17 2 3 1 5 6 7 4 3 2 8 9 3 3 2 3 2 10 
8 1 5 6 7 2 3 4 8 
15 1 5 6 3 2 4 7 8 9 3 2 9 3 2 10 
5 1 5 6 2 3 
3 1 5 6 
28 1 5 6 2 3 7 8 9 9 3 2 2 3 3 2 3 2 3 2 3 2 3 3 2 3 3 2 10 
3 1 5 6 
15 1 5 6 3 4 2 7 8 9 2 3 9 3 2 10 
16 1 5 6 7 2 3 4 8 9 2 3 9 2 3 10 11 
9 1 5 6 2 4 3 7 8 9 
12 1 5 3 4 2 6 8 7 9 9 10 11 
16 1 5 6 3 2 9 2 3 2 2 3 3 2 10 3 2 
29 1 5 6 3 2 4 7 8 12 4 2 4 3 4 3 4 2 4 2 3 9 2 3 9 3 2 3 3 10 
13 1 5 6 2 3 4 7 8 9 9 2 3 10 
21 1 5 6 2 4 3 8 7 9 3 2 3 9 2 2 3 9 3 2 10 11 
12 1 5 6 7 2 3 4 8 9 9 3 10 
29 1 5 6 7 2 4 3 8 9 12 3 4 2 4 2 3 9 3 2 3 4 2 3 4 3 2 2 3 10 
14 1 5 6 7 8 2 3 4 4 9 9 3 2 10 
5 6 1 5 2 3 
10 1 5 6 3 2 9 2 2 9 10 
15 1 5 6 4 3 2 7 8 9 2 3 2 3 2 10 
12 1 5 6 3 4 2 7 8 9 3 2 10 
5 1 5 3 2 6 
11 1 5 6 7 8 2 4 3 9 3 10 
18 1 5 6 2 3 9 2 3 2 2 2 2 2 4 3 2 10 11 
15 1 5 6 3 2 4 8 9 9 2 3 2 3 10 11 
18 1 5 6 2 9 2 2 2 3 2 2 2 2 2 2 3 2 10 
13 1 5 6 7 8 2 4 3 9 2 2 3 10 
16 2 3 1 5 6 4 2 3 7 8 9 2 3 3 2 10 
41 1 5 6 3 2 4 7 8 9 9 12 3 2 4 4 4 2 3 3 4 2 3 2 4 4 3 2 3 2 4 2 4 3 3 2 4 4 2 3 16 11 
6 1 5 6 2 3 2 
6 1 5 6 3 2 4 
9 1 5 6 3 4 2 9 9 10 
13 1 7 6 8 5 4 3 2 9 2 3 10 11 
13 1 5 6 2 3 4 7 8 9 3 2 10 11 
33 1 5 6 4 2 3 9 2 3 2 3 2 3 3 2 2 3 3 2 3 4 3 2 3 3 3 3 2 3 2 3 10 11 
5 1 5 3 2 6 
11 1 5 6 3 4 2 8 9 2 3 10 
8 1 5 6 2 3 4 7 8 
16 1 5 6 4 2 3 9 3 2 3 2 3 2 3 10 11 
14 1 5 6 3 2 4 7 8 9 2 3 3 2 10 
8 1 5 6 4 2 3 7 8 
29 1 5 6 7 8 4 2 3 9 9 2 3 2 2 2 2 2 3 2 2 2 3 2 3 2 2 3 2 15 
10 1 5 6 3 4 2 8 9 7 13 
11 1 5 6 4 2 3 8 9 2 3 10 
20 1 5 6 2 4 3 8 7 9 2 3 9 3 2 9 2 3 2 3 10 
9 1 5 6 8 2 3 4 9 10 
15 1 5 6 7 2 3 8 9 2 2 3 3 2 10 11 
10 1 5 6 3 4 2 7 8 9 10 
13 1 5 6 4 3 2 8 9 3 3 2 10 11 
8 1 5 3 4 2 6 7 8 
12 1 5 6 2 4 3 7 8 9 3 2 10 
17 1 5 6 2 3 4 8 9 9 7 3 2 9 2 3 10 11 
12 1 6 5 7 8 3 2 4 9 9 10 11 
12 1 5 6 7 3 4 2 8 9 3 2 10 
17 1 5 6 3 2 9 2 3 3 2 3 2 2 3 3 2 10 
5 1 5 6 3 2 
13 1 5 6 3 4 2 7 8 9 2 3 10 11 
16 1 5 6 3 2 4 8 7 9 2 3 9 2 3 10 11 
8 1 3 4 2 7 5 6 8 
23 1 5 6 2 3 12 3 2 4 2 2 2 2 4 4 2 3 2 4 2 3 4 13 
5 1 5 6 2 2 
12 1 5 6 2 4 3 8 9 3 2 10 11 
13 1 5 3 4 2 7 6 8 9 3 4 3 10 
3 1 5 6 
5 1 5 6 2 3 
5 1 5 6 3 2 
22 1 5 6 3 2 4 8 7 9 3 2 3 2 3 2 3 2 9 2 3 2 10 
7 1 5 6 3 2 9 10 
13 1 5 6 2 3 4 7 8 9 3 9 3 10 
15 1 5 6 4 3 2 7 8 9 3 2 2 3 10 11 
10 1 5 3 2 6 8 9 4 9 13 
13 1 5 6 7 8 4 2 3 9 2 3 9 10 
12 1 5 6 4 3 2 7 8 9 2 3 10 
14 1 5 6 4 3 2 8 9 9 3 2 3 15 11 
8 1 5 6 3 4 2 7 8 
12 2 1 5 6 3 4 2 8 9 9 2 10 
9 1 5 6 4 3 2 9 10 11 
13 1 5 2 4 3 6 7 8 9 3 2 10 11 
8 1 5 6 7 8 2 4 3 
16 1 5 4 2 3 6 7 8 9 3 2 9 2 3 10 11 
14 1 5 6 4 2 3 7 8 9 9 2 3 10 11 
8 1 5 6 7 2 4 3 8 
15 1 5 3 4 2 6 7 8 9 3 2 2 3 10 11 
6 1 5 6 4 3 2 
11 1 5 6 3 2 4 9 7 8 3 10 
9 1 5 6 4 2 3 9 9 10 
16 1 5 6 7 3 4 2 8 9 2 3 9 3 2 10 11 
18 1 5 6 4 2 3 7 8 9 3 2 9 3 2 2 3 3 10 
21 1 5 6 3 2 4 9 9 3 2 2 3 2 3 2 3 3 2 2 3 14 
14 1 5 6 4 3 2 8 9 7 3 2 3 2 10 
18 1 5 6 7 8 4 3 2 9 9 2 3 3 3 2 3 10 11 
9 1 5 6 3 2 9 3 10 11 
39 1 5 3 2 4 6 7 8 9 12 3 4 2 4 2 3 4 12 4 3 2 4 2 3 2 3 4 9 3 2 3 2 3 2 9 3 2 10 11 
14 1 5 6 4 2 3 7 8 9 3 2 2 3 10 
18 1 5 6 7 8 3 2 4 9 2 2 2 3 9 2 3 3 10 
25 1 5 6 2 3 4 7 8 9 2 3 3 2 2 3 2 9 3 2 2 2 3 3 2 10 
21 1 5 6 2 3 4 7 8 12 4 2 3 4 3 4 2 9 3 2 3 10 
25 2 3 1 5 6 4 2 3 7 8 9 2 3 4 2 3 9 9 3 2 3 2 3 9 13 
23 1 5 3 2 4 6 7 8 12 4 3 2 2 3 4 3 4 2 9 2 3 10 11 
11 1 5 2 3 4 6 8 9 3 2 10 
13 1 5 4 3 2 6 7 8 9 3 2 10 11 
21 1 5 6 7 8 3 4 2 12 2 3 4 4 3 2 4 2 3 9 10 11 
15 1 5 6 2 3 4 7 8 9 3 2 3 2 3 10 
16 1 5 6 2 3 4 7 8 9 9 9 3 2 3 2 10 
12 1 5 6 2 3 4 7 8 9 2 3 10 
10 1 5 6 2 3 4 8 9 4 10 
31 1 5 6 4 3 2 7 8 9 2 3 3 2 9 3 2 3 9 9 3 3 2 3 2 3 3 2 3 3 9 15 
13 1 5 2 3 6 7 8 9 9 3 2 3 10 
14 1 5 3 4 2 6 7 8 9 9 2 3 10 11 
23 1 2 3 4 5 6 8 12 4 2 3 4 2 3 3 2 4 9 2 3 2 3 10 
19 1 5 6 2 3 4 7 8 9 4 3 3 4 2 2 3 2 3 13 
14 1 5 6 2 3 4 8 7 9 2 3 2 3 10 
7 1 5 6 4 3 2 8 
16 1 5 4 3 2 7 6 9 8 3 3 2 3 2 10 11 
15 7 1 5 6 8 2 4 3 9 2 3 2 3 10 11 
16 1 5 6 2 4 3 7 8 9 2 2 3 3 3 10 11 
13 1 5 6 4 3 2 7 8 9 9 3 2 10 
13 1 5 6 4 2 3 7 8 9 2 2 10 11 
12 1 5 6 3 2 9 2 3 9 2 3 10 
16 1 5 6 7 8 4 2 3 9 2 3 9 3 2 3 10 
11 1 5 6 7 2 3 4 8 9 3 2 
13 1 5 6 7 8 3 2 4 9 3 2 10 11 
5 1 5 6 3 2 
13 1 4 2 3 5 6 8 7 9 3 2 10 11 
20 1 5 6 7 2 3 4 8 12 2 3 4 3 4 2 2 4 3 9 13 
17 1 5 6 7 8 2 3 4 9 3 3 2 2 3 3 2 10 
88 2 3 1 5 6 7 4 2 3 8 9 2 3 9 3 2 2 2 3 2 2 2 2 2 3 2 2 2 2 2 2 3 3 2 2 3 2 3 3 2 2 3 2 2 3 2 3 2 3 2 2 2 3 3 2 3 2 2 3 2 12 2 3 4 3 4 2 4 2 3 2 3 4 9 2 2 2 2 3 2 2 3 2 2 3 3 2 15 
10 1 5 6 3 4 2 7 8 9 14 
6 1 5 6 2 3 4 
31 1 5 6 2 3 4 8 7 12 3 4 2 4 4 4 3 4 2 4 4 4 4 4 2 3 9 3 2 2 3 10 
14 1 5 4 2 3 6 7 8 9 3 2 3 2 10 
12 1 5 6 3 4 2 7 8 9 3 2 10 
27 1 5 6 2 3 4 7 8 12 4 2 3 2 3 4 9 2 3 3 2 2 2 3 2 3 10 11 
18 1 5 6 3 4 2 7 8 9 2 3 3 2 2 3 3 3 10 
19 1 5 6 4 3 2 8 7 9 2 3 2 2 3 3 2 2 10 11 
23 1 5 6 4 2 3 7 8 9 3 2 2 3 2 3 2 2 3 2 2 3 10 11 
16 2 3 1 5 6 8 9 2 3 2 3 3 3 2 3 10 
15 1 5 6 7 8 4 2 3 9 3 2 2 3 2 10 
32 1 5 4 3 2 6 7 8 9 3 2 2 3 9 2 3 2 2 3 2 3 2 3 2 3 3 2 3 2 3 14 11 
5 1 5 6 3 2 
18 1 5 6 2 3 4 9 2 3 9 3 2 2 3 2 3 10 11 
20 1 5 4 3 2 6 7 8 9 2 3 3 2 9 2 3 9 2 3 10 
8 2 3 1 5 6 8 9 10 
6 1 5 6 2 4 3 
17 1 5 6 4 3 2 7 8 9 3 2 2 3 3 2 10 11 
11 1 5 6 7 2 3 8 9 3 2 10 
19 1 5 4 2 3 6 7 2 8 9 9 2 3 3 2 2 3 10 11 
11 1 5 6 2 3 8 9 9 9 3 10 
4 1 5 6 2 
11 1 5 6 2 3 4 8 7 9 2 10 
14 1 5 6 7 2 4 3 8 9 9 2 2 3 10 
9 1 5 6 2 4 3 9 7 8 
15 1 5 6 4 2 3 8 9 9 3 2 3 2 10 11 
15 1 5 6 3 4 2 7 8 9 2 3 2 3 10 11 
13 1 5 6 8 2 3 4 7 9 3 2 3 10 
10 1 5 6 4 3 2 7 8 9 10 
5 1 5 2 3 6 
22 1 5 6 4 2 3 8 7 9 2 2 3 2 2 3 2 3 3 2 2 3 10 
29 1 5 6 2 4 3 7 8 9 3 2 2 3 12 2 3 4 4 3 2 4 2 3 9 2 2 3 10 11 
6 1 5 6 3 2 4 
12 1 5 6 3 2 9 2 3 3 2 10 11 
6 1 4 2 3 5 6 
6 1 5 6 3 4 2 
7 1 5 6 2 3 9 10 
16 1 5 2 3 4 6 8 7 9 9 3 2 2 3 10 11 
17 1 5 6 7 8 3 2 4 9 2 3 9 2 3 2 3 10 
7 1 2 4 3 5 6 8 
14 1 5 6 2 3 4 7 8 9 2 3 3 2 10 
9 3 2 1 5 6 9 3 3 10 
14 1 5 6 3 4 2 7 8 9 2 2 3 10 11 
18 1 5 4 3 2 6 7 8 9 2 3 4 3 2 2 3 10 11 
13 1 5 6 7 8 2 4 3 9 2 3 10 11 
5 1 5 6 2 3 
9 1 5 2 3 6 7 8 13 9 
15 1 5 6 4 2 3 8 9 3 2 9 2 3 3 10 
8 1 5 3 4 2 6 7 8 
29 1 5 6 4 2 3 7 8 12 2 4 3 2 3 4 4 4 3 2 9 2 3 2 3 3 2 3 10 11 
16 1 6 5 8 2 3 7 9 3 2 3 2 3 3 2 10 
13 1 5 6 8 2 4 3 7 9 2 3 9 14 
15 2 3 1 5 6 9 3 2 9 3 2 3 2 3 14 
37 1 6 5 3 2 4 4 7 8 12 4 2 3 4 3 4 2 9 2 3 2 2 3 2 3 2 3 2 3 2 3 2 2 3 2 3 10 
13 1 5 6 4 3 2 9 9 2 3 3 2 16 
170 1 5 6 7 4 3 2 8 9 2 3 12 3 2 4 2 2 4 2 3 4 3 2 4 3 4 2 3 4 2 4 2 3 3 2 4 3 2 4 4 2 3 4 3 2 2 3 4 3 2 4 3 2 4 4 2 3 4 3 2 4 2 3 2 3 2 4 2 4 3 4 2 3 3 4 2 3 2 4 3 4 2 12 3 4 2 2 2 3 4 4 3 4 2 3 2 4 3 4 2 3 4 2 4 3 2 4 2 3 3 2 4 2 3 4 3 2 4 4 2 3 4 2 3 4 2 3 4 3 2 4 3 2 2 3 4 4 2 3 3 4 2 2 3 4 4 3 2 3 4 2 3 4 2 2 4 3 2 4 3 3 4 2 2 9 2 3 2 10 11 
35 1 5 6 7 4 2 3 8 12 3 2 4 2 4 3 3 2 4 4 3 2 9 2 3 3 2 3 2 3 2 2 3 3 2 10 
20 1 5 6 3 2 9 3 2 3 2 2 2 2 2 2 2 2 2 3 10 
15 1 5 6 4 2 3 7 8 9 9 3 3 3 10 11 
19 1 5 6 3 2 4 7 8 9 2 4 3 9 3 2 2 3 10 11 
8 1 5 4 3 2 6 7 8 
12 1 5 6 4 3 2 7 8 9 2 3 10 
7 1 5 3 2 6 9 10 
40 1 5 6 2 4 3 8 7 12 3 4 2 4 2 4 3 2 4 4 2 3 4 9 2 3 3 3 3 2 3 2 3 2 3 2 3 2 9 10 11 
7 1 5 6 2 3 8 7 
9 1 5 7 2 3 2 4 6 8 
15 1 5 6 2 3 7 8 9 3 2 3 2 3 2 10 
16 1 5 6 7 3 4 2 8 9 2 3 2 3 2 10 11 
18 1 5 6 3 4 2 7 8 9 9 3 2 3 2 3 2 10 11 
13 1 7 5 6 4 2 3 8 9 2 3 10 11 
28 1 5 6 4 3 2 7 8 9 3 2 3 9 3 2 3 3 2 2 2 3 3 2 3 3 2 2 10 
8 1 5 6 3 2 4 8 7 
26 1 5 6 3 4 2 7 8 9 2 3 3 2 3 2 2 3 3 2 2 3 3 2 3 3 10 
11 1 5 6 2 3 4 8 7 9 9 13 
5 1 5 6 3 2 
8 1 5 6 3 4 2 7 8 
23 1 7 5 6 3 4 2 8 9 2 9 4 3 2 4 2 3 2 3 4 3 2 13 
41 1 5 6 4 2 3 7 8 9 2 3 9 2 3 4 3 2 9 2 12 3 4 2 2 2 3 4 2 9 2 3 2 2 2 2 3 2 3 2 15 11 
18 1 5 6 7 2 3 4 8 9 9 3 2 2 3 3 2 10 11 
11 1 5 6 4 3 2 7 8 9 2 3 
12 1 5 3 4 2 6 7 8 9 3 2 10 
14 1 7 5 6 3 4 2 8 9 9 2 3 9 10 
15 1 5 6 7 8 2 3 4 9 3 2 2 3 10 11 
33 3 2 1 5 6 9 3 2 12 2 3 4 2 2 12 2 3 4 2 2 2 4 3 2 4 2 3 3 4 2 9 10 11 
13 1 5 6 8 3 2 9 2 3 7 3 2 10 
15 1 5 4 2 3 6 7 8 9 2 3 9 3 2 10 
6 2 1 5 6 2 3 
16 1 5 6 7 8 2 3 4 9 3 2 9 2 3 2 10 
20 1 5 2 4 3 6 7 8 9 3 2 2 3 2 3 3 2 3 2 13 
8 1 5 6 2 3 4 7 8 
27 1 5 6 4 2 3 9 9 8 7 3 2 3 2 3 3 2 9 12 4 2 3 3 2 4 9 10 
5 1 5 6 2 3 
28 1 5 6 4 2 3 8 7 9 12 4 3 2 3 2 4 3 2 4 9 3 2 3 2 3 2 10 11 
23 1 5 6 2 4 3 7 8 9 2 3 3 2 2 2 3 2 3 2 2 3 15 11 
16 1 2 3 4 5 6 7 8 9 9 3 2 3 2 10 11 
7 3 2 1 2 3 5 6 
5 1 5 6 2 3 
7 1 5 6 2 9 10 11 
6 1 5 6 4 2 3 
8 1 3 2 5 6 8 9 10 
16 1 5 7 2 3 4 6 8 9 2 3 9 3 2 10 11 
15 1 5 6 4 2 3 7 8 9 2 3 2 3 10 11 
28 1 2 3 4 5 6 8 7 9 12 4 3 2 4 3 2 2 3 4 3 2 4 3 4 2 9 3 10 
20 1 5 6 2 3 4 7 8 9 12 3 4 2 3 4 2 9 3 2 10 
25 1 5 6 2 3 4 7 8 9 3 2 4 3 2 3 2 2 3 2 3 2 3 2 3 10 
17 1 5 6 7 4 2 3 8 9 9 3 2 3 2 3 10 11 
12 1 5 6 7 2 3 4 8 9 9 10 11 
16 1 5 6 7 2 3 8 9 3 2 3 2 2 3 10 11 
8 1 5 6 2 3 4 7 8 
10 1 5 2 3 4 7 9 6 8 10 
13 1 5 6 7 4 3 2 8 9 9 2 3 10 
11 1 5 6 2 3 4 8 9 2 3 10 
13 1 5 6 2 4 3 8 9 2 3 3 2 10 
13 1 5 6 7 2 4 3 8 9 2 3 10 11 
17 1 6 5 3 2 7 8 4 12 2 3 2 4 2 3 4 2 
16 1 5 2 3 4 6 7 8 9 2 3 3 3 2 10 11 
34 1 5 6 4 2 3 7 8 12 4 4 2 4 3 4 2 4 4 2 3 4 4 3 4 2 2 3 4 2 3 4 9 10 11 
7 1 5 6 4 2 3 9 
22 1 5 6 7 3 2 4 8 9 3 2 2 2 3 4 4 2 3 3 2 10 11 
18 7 1 5 6 2 3 4 8 9 2 3 4 3 2 3 2 10 11 
9 1 5 6 8 4 2 3 9 13 
27 1 5 6 2 3 4 7 8 9 9 3 2 4 2 2 3 3 2 2 3 2 3 3 2 2 3 10 
12 1 5 6 7 8 3 4 2 9 3 2 10 
11 1 5 6 7 3 2 4 8 9 3 2 
22 1 5 6 9 12 2 3 4 2 4 3 2 3 4 9 3 2 2 3 3 2 10 
15 1 5 6 7 8 2 4 3 9 9 2 3 3 2 14 
14 1 5 2 3 6 7 4 8 9 3 2 3 2 10 
8 1 5 6 7 3 4 2 8 
6 1 5 6 3 2 8 
10 1 5 3 2 4 9 6 7 8 10 
11 1 5 6 4 2 3 9 9 3 2 10 
16 1 5 6 3 2 7 8 9 2 3 9 3 2 3 10 11 
5 1 5 6 2 3 
10 1 7 5 4 2 3 6 8 9 10 
19 1 6 5 7 4 3 2 8 9 3 4 2 3 2 3 2 2 3 13 
22 1 5 6 7 3 2 4 8 9 4 3 2 3 2 4 3 2 4 2 3 10 11 
16 1 5 6 2 4 3 7 8 9 2 3 3 2 3 10 11 
8 1 5 6 3 4 2 7 8 
5 1 5 6 2 3 
17 1 5 6 4 2 3 7 8 9 3 2 9 2 3 3 2 10 
14 1 5 2 3 6 9 2 3 2 2 3 3 2 10 
3 1 5 6 
15 1 5 6 2 3 4 7 8 9 2 3 9 2 3 10 
11 1 5 6 4 3 2 7 8 9 9 10 
15 1 5 4 3 2 6 7 8 9 9 3 2 2 3 13 
16 1 5 6 2 3 4 7 8 12 2 3 4 9 2 3 10 
13 1 5 6 4 2 3 7 8 9 2 9 2 10 
30 1 5 6 3 2 4 7 8 9 3 2 2 3 9 9 2 3 2 3 2 2 3 3 2 2 3 2 2 3 13 
12 1 7 6 8 5 4 2 3 9 2 3 10 
14 1 5 6 2 3 4 7 8 9 3 2 3 2 10 
12 1 5 6 3 2 4 7 8 9 3 2 10 
13 1 6 8 5 3 2 4 7 9 3 2 9 10 
8 1 5 6 3 4 2 7 8 
30 1 5 6 2 3 4 7 8 9 9 3 2 2 3 2 2 3 3 2 3 2 2 2 3 2 3 3 2 10 11 
8 1 5 3 2 4 6 9 13 
10 1 5 6 2 4 3 8 9 3 10 
13 1 5 6 2 3 4 7 8 9 9 2 3 10 
13 1 5 6 2 3 4 7 8 9 2 3 10 11 
18 1 5 3 2 4 6 7 8 9 2 2 2 3 3 2 2 3 13 
11 1 5 3 2 6 9 3 2 3 10 11 
21 1 5 6 4 2 3 7 8 9 4 3 2 9 3 4 2 2 3 3 10 11 
16 1 5 6 4 3 2 8 9 3 2 9 3 3 2 10 11 
5 1 5 6 3 2 
12 1 5 6 8 2 4 3 9 3 3 2 10 
5 1 5 6 9 10 
10 1 5 6 4 2 3 8 9 3 10 
8 1 5 6 7 8 3 4 2 
12 1 5 6 2 3 12 2 2 2 3 3 13 
15 1 5 6 7 4 2 3 8 9 2 3 2 3 10 11 
12 1 5 6 4 2 3 9 9 3 2 10 11 
12 1 5 6 3 2 4 7 8 9 3 2 15 
13 1 5 6 4 2 3 7 8 9 2 3 10 11 
14 1 5 6 2 3 4 7 8 9 9 2 3 10 11 
12 1 5 6 2 4 3 7 8 9 3 2 10 
21 1 5 6 2 4 3 7 8 9 2 3 3 3 2 2 3 10 11 3 4 2 
23 1 5 6 2 4 3 7 8 9 3 2 3 2 3 2 2 3 2 3 2 3 10 11 
11 1 5 6 7 8 3 2 4 9 10 11 
17 1 5 6 4 3 2 7 8 9 2 3 3 2 2 3 10 11 
15 1 5 6 2 3 4 7 8 9 2 3 9 2 3 10 
8 1 5 6 2 4 3 7 8 
9 1 5 6 3 4 2 7 8 9 
5 1 5 6 2 3 
10 1 5 6 4 3 2 8 7 9 10 
9 1 5 6 3 2 4 7 8 5 
16 1 5 6 4 2 3 7 8 9 3 3 2 3 2 10 11 
9 1 5 6 2 4 3 7 8 9 
12 1 5 6 2 3 4 8 7 9 3 2 10 
12 1 5 6 2 4 3 8 7 9 9 9 10 
19 1 5 6 7 8 2 3 4 9 3 2 3 2 9 3 2 3 2 13 
22 1 5 6 3 2 4 7 8 12 3 4 2 4 4 3 2 9 3 2 3 10 11 
14 1 5 2 3 9 6 9 2 3 2 3 2 3 14 
5 1 5 6 3 2 
11 7 1 5 6 2 3 4 8 9 10 11 
13 1 5 6 7 3 4 2 8 9 3 2 3 10 
8 1 5 6 2 3 4 9 13 
15 1 5 6 2 3 4 7 8 9 3 2 9 2 3 14 
16 5 1 6 7 8 2 3 4 9 9 3 2 3 2 14 11 
18 3 4 2 1 5 6 7 8 9 2 3 3 2 3 2 2 3 14 
6 1 3 2 5 6 8 
17 1 5 6 7 8 4 2 3 9 4 2 3 3 2 2 3 10 
13 1 5 6 2 3 4 7 8 9 2 3 3 10 
22 1 5 6 3 4 2 7 8 2 3 4 12 2 4 2 4 2 3 4 3 2 13 
13 1 5 6 7 3 4 2 8 9 3 3 3 14 
7 1 5 6 2 4 3 8 
15 7 1 5 6 8 3 2 4 9 9 2 3 2 3 10 
48 1 5 6 3 4 2 7 8 9 9 9 2 2 3 2 3 12 2 3 4 2 2 2 2 2 2 2 3 4 2 2 2 2 2 2 2 2 4 3 4 2 3 9 2 2 2 10 11 
6 1 5 6 2 3 4 
16 1 5 6 2 3 9 3 2 9 3 2 2 3 3 2 13 
45 1 5 6 4 3 2 7 8 3 4 2 12 4 2 3 2 3 4 2 3 4 4 2 3 3 4 2 2 3 4 2 3 4 9 2 2 3 2 2 3 2 2 3 15 11 
23 1 5 6 3 2 4 7 8 9 3 3 2 3 2 2 3 2 3 3 2 3 2 10 
39 1 5 2 3 6 7 8 9 2 3 2 3 3 2 3 3 2 3 2 3 2 3 2 2 3 3 2 2 3 3 3 3 2 3 2 3 3 2 10 
22 1 5 6 7 4 2 3 8 9 9 4 2 3 2 3 2 3 3 2 3 10 11 
15 1 5 6 3 4 2 7 8 9 2 3 2 2 10 11 
15 7 1 5 6 8 4 2 3 9 9 3 2 2 10 11 
6 1 5 6 2 3 4 
12 1 5 6 4 2 3 7 8 9 3 10 11 
10 1 5 6 2 3 4 7 8 9 10 
12 1 5 6 2 4 3 7 8 9 3 2 10 
10 1 5 6 2 3 4 7 8 9 10 
13 1 5 6 3 2 4 7 8 9 2 3 10 11 
20 1 5 6 2 4 3 7 8 9 3 2 2 3 2 3 3 2 3 2 14 
15 1 5 6 2 4 3 7 8 9 2 3 9 3 2 10 
16 1 5 6 7 8 2 3 4 9 9 3 2 3 2 2 10 
6 1 5 6 2 3 4 
21 1 5 6 7 4 2 3 8 9 2 3 2 3 3 2 2 3 2 3 14 11 
23 1 5 6 3 2 4 7 8 12 4 4 3 2 9 2 3 2 3 2 3 2 10 11 
14 1 5 6 2 3 4 7 4 2 3 8 9 10 11 
8 1 5 6 3 4 2 7 8 
13 1 5 6 7 2 3 4 8 9 2 3 10 11 
12 1 5 6 4 3 2 8 9 7 3 2 10 
9 1 5 6 2 3 4 9 9 10 
10 1 5 6 4 3 2 7 8 9 10 
37 1 5 6 4 2 3 8 12 4 2 3 2 3 4 2 3 4 3 2 4 3 2 4 4 2 3 2 3 4 9 3 2 3 2 2 9 10 
22 1 5 6 4 3 2 9 2 3 9 2 3 2 3 2 3 2 3 2 3 10 11 
14 1 5 6 2 3 4 7 8 9 2 3 3 2 10 
16 1 5 6 4 3 2 7 8 9 9 3 2 3 2 10 11 
14 1 5 6 3 2 4 8 9 9 2 3 2 3 10 
13 1 5 6 7 4 2 3 8 9 9 2 3 10 
29 1 2 3 4 5 6 8 9 9 2 3 9 12 4 3 2 4 3 2 2 4 3 9 2 3 3 2 3 10 
12 1 5 7 2 3 4 6 8 9 3 10 11 
17 1 5 6 7 8 2 4 3 9 9 2 3 3 2 3 2 10 
16 1 5 6 4 2 3 7 8 9 9 2 3 2 3 10 11 
13 1 5 3 4 2 6 7 8 9 3 2 9 10 
11 1 5 6 2 3 4 7 8 9 2 3 
11 1 5 6 7 2 4 3 8 9 10 11 
17 1 5 6 7 4 3 2 8 9 3 4 2 9 2 3 10 11 
5 1 5 6 2 3 
12 1 2 3 4 5 6 8 7 9 2 3 10 
16 1 5 6 2 3 4 7 8 9 2 3 9 2 3 9 10 
18 1 5 3 4 2 6 7 8 9 2 3 2 2 3 2 9 10 11 
18 1 5 3 2 4 6 7 8 9 2 3 2 3 2 3 2 10 11 
17 1 5 4 3 2 7 6 8 9 9 3 2 3 2 3 10 11 
13 1 5 6 3 2 4 7 8 9 2 3 2 15 
12 1 5 6 7 8 4 2 3 9 2 3 10 
14 1 5 6 7 8 2 4 3 9 3 2 3 2 10 
11 1 5 6 3 2 4 9 3 2 10 11 
9 1 5 6 7 2 4 3 8 9 
14 1 5 6 4 2 3 8 7 9 3 2 2 10 11 
12 1 5 6 3 4 2 9 2 3 2 3 10 
15 1 5 6 2 3 7 8 9 2 2 2 2 2 10 11 
3 1 5 6 
15 1 5 6 8 7 4 3 2 9 9 2 3 2 3 10 
16 1 2 4 3 5 6 7 8 9 9 3 3 2 3 2 10 
8 1 5 6 3 4 2 7 8 
13 1 5 6 2 3 4 8 9 2 3 7 10 11 
14 1 5 6 7 8 3 4 2 9 2 3 3 2 10 
20 1 5 6 7 4 3 2 8 9 3 2 9 3 2 3 2 3 2 3 10 
14 1 2 4 3 5 6 7 8 9 9 3 2 10 11 
38 1 5 2 3 4 6 7 8 9 9 2 3 2 2 3 2 3 2 3 3 2 3 2 3 3 2 3 3 3 2 3 3 2 2 2 2 3 13 
19 1 5 6 7 4 3 2 8 9 9 2 3 4 2 3 3 2 10 11 
34 2 3 1 5 6 8 9 3 2 9 3 2 9 12 2 4 3 3 4 2 2 2 4 3 9 2 3 2 3 2 3 3 2 10 
9 1 5 6 7 2 4 3 8 9 
20 1 5 2 4 3 6 9 9 3 2 2 3 3 2 3 3 2 3 3 15 
6 1 5 6 2 9 10 
14 1 5 6 4 2 3 7 8 9 2 3 3 2 10 
17 1 5 6 4 2 3 7 8 9 4 9 4 2 3 4 3 10 
8 1 5 6 4 2 3 8 7 
3 1 5 6 
10 1 5 6 3 4 2 7 8 9 10 
10 1 4 3 2 5 6 7 8 9 10 
16 1 5 6 3 4 2 7 8 9 3 2 4 9 3 2 10 
12 1 5 6 2 4 3 7 8 9 2 3 10 
8 1 5 6 3 4 2 7 8 
10 1 5 6 4 3 2 8 2 3 7 
8 1 5 6 7 8 4 2 3 
14 1 5 6 7 8 4 2 3 9 2 3 2 3 13 
16 1 3 2 4 5 6 7 8 9 3 2 3 2 2 3 10 
8 1 5 3 2 6 7 4 8 
15 1 5 6 7 8 2 4 3 9 3 4 2 2 3 10 
8 1 5 2 3 6 9 10 11 
19 1 5 6 2 3 9 2 3 2 3 3 2 3 2 2 3 3 2 15 
16 1 5 2 3 4 6 7 8 9 3 2 9 3 2 3 10 
11 1 7 5 6 8 4 3 2 9 3 10 
9 1 5 2 3 4 6 8 9 7 
14 1 5 6 2 3 4 7 8 9 9 2 3 10 11 
9 1 5 6 3 2 4 7 8 9 
3 1 5 6 
10 1 5 6 2 4 3 7 8 9 13 
17 1 5 6 2 3 4 7 8 9 3 2 2 3 2 3 10 11 
15 1 5 6 4 2 3 7 8 9 3 2 2 3 10 11 
5 1 5 6 3 2 
14 1 5 6 4 3 2 7 8 9 3 2 3 2 10 
8 1 5 2 4 3 6 7 8 
21 1 5 6 7 8 2 4 3 9 2 3 3 2 3 2 3 2 3 2 10 11 
12 1 5 6 4 2 3 7 8 9 2 3 10 
7 1 5 6 3 2 4 8 
21 1 7 5 2 3 4 6 8 9 4 2 9 9 2 3 3 2 2 3 2 10 
15 1 3 4 2 5 6 7 8 9 9 2 3 3 2 10 
13 1 5 4 2 3 6 7 8 9 2 3 9 10 
23 1 5 6 4 2 3 7 8 9 2 3 9 2 3 2 3 2 3 2 3 2 3 10 
20 1 5 2 4 3 6 7 8 9 3 2 2 3 2 3 9 3 2 10 11 
11 6 7 8 1 5 4 3 2 4 3 2 
6 1 5 6 2 3 5 
13 2 1 5 6 7 3 2 4 8 9 3 2 10 
16 1 5 6 4 2 3 7 8 9 9 2 3 3 2 10 11 
13 1 5 6 4 2 3 7 8 9 9 3 10 11 
15 2 3 1 5 6 7 4 8 9 9 3 2 3 3 10 
30 1 5 6 4 3 2 7 8 9 4 2 3 2 3 3 2 3 2 3 2 3 3 2 2 3 2 3 9 9 13 
18 1 5 6 4 3 2 7 8 9 9 4 3 2 2 3 2 3 10 
16 1 5 6 3 2 4 7 8 9 3 2 3 2 3 2 10 
12 1 5 6 3 2 4 7 8 9 3 3 10 
14 1 5 6 4 3 2 8 7 9 9 2 3 10 11 
15 1 5 6 3 4 2 7 8 9 2 3 9 3 2 10 
19 1 5 6 7 8 2 3 4 9 4 2 3 9 9 2 3 2 3 10 
22 1 5 6 3 2 4 7 8 9 4 3 2 2 3 2 2 2 2 2 9 10 11 
14 2 1 5 6 7 2 3 4 8 9 2 3 10 11 
14 5 1 6 3 2 4 7 8 9 2 3 9 10 11 
18 1 5 6 7 2 3 4 8 12 3 4 2 12 9 3 2 10 11 
16 1 5 6 3 4 2 7 8 9 3 2 2 3 2 3 10 
10 1 5 6 2 3 9 3 2 3 10 
13 1 5 6 7 2 4 3 8 9 9 3 2 10 
6 1 5 6 2 3 4 
17 1 5 3 2 4 6 7 8 9 3 2 2 3 3 2 10 11 
14 1 5 6 4 3 2 8 9 3 2 9 2 3 10 
13 2 3 1 5 2 3 4 6 7 8 9 3 10 
24 1 5 6 2 4 3 8 7 9 9 2 3 3 2 3 9 9 3 9 2 3 3 2 10 
17 1 5 6 4 3 2 8 9 3 2 9 3 2 2 3 10 11 
15 6 1 5 3 2 4 8 7 9 2 3 9 2 3 13 
10 1 5 6 7 4 2 3 8 9 10 
8 1 5 6 2 4 3 7 8 
17 1 7 5 6 4 2 3 8 12 4 2 4 3 9 3 2 10 
30 5 2 3 4 2 1 12 4 2 3 3 4 2 3 2 4 2 4 3 2 3 4 4 3 2 9 2 3 10 11 
13 2 1 5 6 3 4 2 7 8 9 3 2 10 
12 1 5 6 2 3 4 7 8 9 2 3 10 
12 1 5 6 4 3 2 8 9 3 3 2 10 
14 1 5 6 3 4 2 8 7 9 3 2 3 10 11 
5 1 5 6 2 3 
29 1 5 6 7 3 2 4 8 9 3 2 2 3 9 9 9 3 2 9 2 2 3 3 2 2 3 2 3 13 
5 1 5 6 3 2 
20 1 5 6 2 4 3 7 8 9 2 3 4 3 2 9 3 2 2 3 10 
15 1 5 6 7 8 2 3 4 9 3 2 2 3 10 11 
8 1 5 6 3 4 2 7 8 
5 1 5 6 3 2 
8 1 5 6 2 4 3 8 7 
12 3 2 1 5 6 4 3 2 7 8 9 13 
84 1 5 6 7 8 3 2 4 9 12 4 2 3 4 2 3 4 4 2 3 4 2 3 4 2 3 4 2 3 2 3 4 4 2 3 2 3 4 2 3 4 4 2 3 3 4 2 2 3 4 3 2 4 3 4 2 2 3 4 2 3 4 4 2 3 3 4 2 2 3 4 2 3 4 3 4 2 2 4 3 4 9 9 10 
10 1 5 6 4 2 3 7 8 9 10 
22 1 5 3 2 4 6 9 2 3 2 3 3 2 3 2 2 3 3 2 2 3 13 
6 1 5 6 2 3 4 
33 1 5 6 2 3 4 7 8 9 9 3 2 12 3 4 2 2 4 3 9 3 2 9 3 2 2 3 3 2 3 2 3 16 
14 1 5 6 2 4 3 7 8 9 2 9 3 2 10 
12 1 5 6 2 3 8 7 9 2 2 2 13 
17 1 5 4 2 3 6 7 8 9 9 3 2 2 3 3 10 11 
13 1 5 4 3 2 6 7 8 9 9 2 3 10 
15 1 5 6 3 2 4 8 9 7 3 2 3 2 10 11 
18 1 5 7 6 4 3 2 8 9 9 2 3 2 3 2 3 10 11 
18 1 5 3 4 2 6 7 8 9 3 2 3 2 2 2 3 10 11 
5 1 5 6 3 2 
3 1 5 6 
6 1 5 6 3 4 2 
8 1 5 6 4 2 3 7 8 
16 1 5 6 2 3 9 3 3 2 3 2 2 3 2 3 10 
8 1 5 6 3 4 2 7 8 
12 1 4 2 3 5 6 9 2 3 3 2 10 
23 3 1 5 6 7 4 2 3 8 9 12 2 4 3 4 3 2 9 2 3 2 3 10 
14 1 5 6 7 8 4 2 3 9 3 2 9 10 11 
3 1 5 6 
9 1 2 3 4 5 6 7 8 9 
17 1 5 4 2 3 6 8 7 9 9 3 2 2 3 3 2 10 
3 1 5 6 
13 1 5 6 3 4 2 8 9 7 2 3 10 11 
21 1 5 6 2 3 4 7 8 9 4 9 9 9 3 2 3 2 3 2 9 10 
8 1 5 6 2 3 4 7 8 
15 1 5 6 2 3 4 7 8 9 2 3 9 3 2 10 
24 1 5 6 4 3 2 8 9 2 3 9 2 3 2 3 2 3 3 2 3 2 2 3 10 
40 1 5 6 2 3 4 4 7 8 3 2 4 12 4 2 3 4 4 4 2 3 9 2 3 4 3 2 2 3 4 9 2 3 2 3 2 3 3 2 13 
32 1 5 6 3 2 7 8 12 4 4 2 4 3 4 4 4 2 3 4 2 3 9 2 3 3 2 3 2 3 2 3 10 
6 1 5 6 2 3 4 
18 1 5 6 3 4 2 7 8 9 9 2 3 2 3 2 2 10 11 
5 1 5 6 2 3 
22 1 5 3 4 2 7 9 6 8 12 3 4 2 2 3 4 9 2 3 3 2 10 
7 1 5 6 3 2 9 10 
10 1 5 6 2 3 4 7 8 3 2 
17 1 7 5 6 4 2 3 8 9 3 3 2 9 9 2 3 10 
21 6 8 7 1 5 3 2 4 9 9 3 2 9 2 3 2 9 2 2 10 11 
14 1 5 6 2 3 4 8 9 3 2 2 3 10 11 
61 1 5 6 2 3 4 7 8 9 12 2 3 4 4 2 3 2 3 4 3 4 2 3 4 2 2 3 4 3 4 2 4 3 2 3 4 2 4 2 3 4 2 3 3 2 4 4 3 2 2 3 4 9 3 2 9 9 2 9 10 11 
10 1 5 6 2 3 4 7 8 2 3 
15 1 5 3 2 4 6 8 9 9 2 3 2 3 15 11 
10 1 5 6 4 3 2 8 9 2 10 
14 1 5 6 2 3 7 8 9 2 3 9 3 3 10 
8 1 2 4 3 5 6 8 7 
8 1 5 6 3 2 7 8 4 
12 1 5 6 3 4 2 7 8 9 2 3 13 
6 1 5 6 2 2 3 
24 1 5 6 3 2 4 7 8 9 3 2 4 2 3 2 3 2 3 3 2 3 2 14 11 
16 7 1 5 6 4 2 3 8 9 2 3 4 3 4 2 13 
15 1 7 5 2 3 4 6 8 9 9 2 3 3 10 11 
14 1 5 6 4 2 3 7 8 9 3 2 2 3 10 
11 1 5 6 7 2 3 4 8 9 10 11 
12 1 5 6 2 3 4 7 8 9 3 2 10 
8 1 7 5 6 4 3 2 8 
16 1 5 2 3 4 6 7 8 9 2 3 2 3 2 3 10 
15 1 5 6 3 4 2 9 2 3 2 9 4 3 2 13 
17 1 5 6 2 3 4 8 9 2 3 4 9 7 3 2 10 11 
16 1 5 6 7 4 3 2 8 9 2 3 2 3 2 3 10 
21 1 5 6 4 2 3 8 12 3 2 4 2 3 4 9 9 2 3 3 2 10 
9 1 5 6 4 3 2 9 10 11 
23 1 5 6 2 3 9 2 9 2 2 2 2 2 2 2 2 3 2 2 2 2 2 16 
5 1 5 6 9 10 
8 1 5 6 4 2 3 7 8 
14 1 5 6 4 2 3 9 3 2 3 2 2 3 10 
3 1 5 6 
37 1 5 6 2 3 4 8 9 3 2 12 2 3 4 2 3 4 4 3 2 2 3 4 3 4 2 4 3 2 4 2 3 2 4 3 9 10 
8 1 5 6 2 3 4 7 8 
14 1 5 6 2 4 3 7 8 9 3 2 3 2 14 
17 1 5 6 3 2 4 7 8 12 3 2 4 9 9 2 3 15 
11 1 5 6 3 2 9 3 2 2 3 16 
18 1 5 6 4 2 3 7 8 9 2 3 2 3 2 3 2 3 10 
5 1 5 6 3 2 
20 1 5 6 7 8 3 2 4 12 3 4 2 4 3 2 9 3 2 10 11 
12 1 7 5 6 4 2 3 8 9 3 2 10 
13 1 6 7 8 5 2 4 3 9 9 2 3 10 
12 1 5 6 2 3 4 7 8 9 2 3 10 
15 1 5 6 3 4 2 7 8 9 9 3 2 3 3 10 
17 1 5 6 7 4 2 3 8 9 2 3 2 2 3 3 2 10 
14 1 5 6 3 4 2 7 8 9 9 2 3 3 10 
21 1 5 6 2 4 3 7 8 9 3 2 4 4 3 9 3 4 2 3 9 10 
14 1 5 4 2 3 6 7 8 9 2 3 9 3 10 
12 1 5 6 4 3 2 7 8 9 3 3 10 
10 1 5 6 2 3 9 2 3 10 11 
11 1 5 6 2 4 3 7 8 9 10 11 
15 1 5 6 3 4 2 7 8 9 3 2 2 3 14 11 
12 1 5 6 7 2 3 4 8 9 3 3 10 
8 1 5 2 3 4 6 7 8 
15 1 5 6 7 3 2 4 8 9 9 2 3 3 2 10 
19 1 5 6 7 3 2 4 8 9 2 3 9 2 3 3 2 3 2 14 
11 1 5 6 7 8 2 3 4 9 3 10 
5 1 5 6 2 3 
13 1 5 6 3 4 2 9 3 2 4 2 3 10 
11 1 5 6 7 8 3 2 4 12 4 13 
33 1 5 6 7 8 4 2 3 12 2 3 4 3 4 2 4 3 2 4 9 3 2 2 3 3 2 3 2 3 2 2 3 10 
13 1 5 6 3 2 4 8 9 2 3 2 3 10 
14 1 5 6 2 4 3 7 8 9 4 9 2 3 10 
12 1 5 6 2 4 3 7 8 9 3 2 10 
15 1 5 6 7 2 4 3 8 9 3 2 3 2 10 11 
5 1 5 2 3 6 
12 1 5 6 3 4 2 9 9 3 3 3 10 
27 1 5 6 2 4 3 9 9 12 4 2 3 2 4 7 8 2 3 4 4 2 3 9 2 2 10 11 
14 1 5 6 3 2 4 7 8 9 2 3 2 3 10 
11 1 5 4 2 3 6 7 8 9 3 10 
8 1 5 6 3 4 2 7 8 
19 1 5 6 7 2 4 3 8 9 3 2 4 4 3 2 2 3 4 16 
8 1 5 6 3 2 4 7 8 
13 1 5 6 4 2 3 7 8 9 2 3 10 11 
19 1 5 2 4 3 12 6 7 8 2 4 3 3 4 2 9 2 3 10 
15 1 5 6 4 3 2 7 8 9 2 3 2 3 10 11 
14 1 5 6 3 4 2 7 8 9 3 2 2 10 11 
8 1 5 6 7 3 2 4 8 
5 1 5 6 3 2 
18 1 5 6 3 2 4 7 8 9 3 2 3 2 3 3 2 15 11 
11 1 7 5 6 3 2 8 9 2 3 10 
8 1 5 6 7 2 3 4 8 
5 1 5 6 2 3 
17 7 1 5 6 8 2 3 4 9 9 3 2 3 2 3 10 11 
5 1 5 6 2 3 
10 1 5 6 2 3 4 9 2 3 4 
15 1 5 6 3 2 4 7 8 9 2 3 9 3 2 10 
15 1 5 6 3 2 4 7 8 9 4 9 2 3 10 11 
17 1 7 5 6 2 3 4 8 12 2 3 4 9 2 9 10 11 
21 1 5 6 3 4 2 7 8 9 2 3 2 3 3 2 3 2 3 2 10 11 
5 1 5 6 2 3 
15 1 5 6 4 3 2 7 8 9 3 2 3 2 10 11 
20 1 5 6 7 8 3 4 2 12 2 3 4 4 3 2 9 3 3 2 10 
35 1 5 6 4 2 3 7 8 9 9 3 2 3 12 4 3 2 4 9 9 3 2 3 2 3 2 3 2 3 2 3 2 3 10 11 
11 1 5 6 3 2 4 8 7 9 2 3 
9 1 5 6 7 3 2 4 8 4 
24 1 5 6 4 2 3 8 9 3 2 3 2 3 2 3 2 3 3 2 10 11 3 2 4 
12 1 5 6 2 3 4 7 8 9 9 2 10 
3 1 5 6 
17 1 5 6 7 8 3 2 4 9 3 2 3 2 2 3 3 10 
12 1 5 6 2 3 4 7 8 9 3 10 11 
18 1 5 6 3 4 2 8 9 2 3 9 7 3 2 2 3 10 11 
9 1 5 6 2 3 9 9 10 11 
12 1 5 6 7 8 4 2 3 9 3 10 11 
13 1 5 6 2 3 4 7 8 9 9 2 10 11 
8 1 5 2 3 4 6 7 8 
3 1 5 6 
15 1 5 6 8 3 4 2 7 9 3 2 9 3 2 10 
12 7 1 5 2 3 4 6 8 12 4 3 2 
15 1 5 6 7 4 2 3 8 12 4 3 2 9 9 10 
23 1 5 6 7 8 3 2 4 9 2 3 2 3 2 3 9 2 3 3 2 2 3 15 
16 1 5 6 2 3 4 7 8 9 9 3 2 4 2 3 10 
9 1 5 6 2 3 9 2 10 11 
8 1 5 6 7 3 2 4 8 
14 1 5 6 3 2 4 7 8 9 2 3 2 3 10 
10 1 5 6 7 8 2 3 4 9 10 
30 2 3 1 5 6 3 4 2 7 8 9 2 3 9 3 2 2 2 3 2 3 3 2 3 2 2 3 2 3 10 
13 1 5 6 7 2 3 4 8 9 2 3 10 11 
31 7 1 5 6 4 2 3 8 12 2 3 4 3 4 2 9 2 3 2 3 2 3 2 3 3 2 2 3 2 3 10 
6 1 5 6 4 2 3 
13 1 5 6 7 8 2 4 3 9 2 3 10 11 
18 1 5 6 7 4 2 3 8 12 3 2 4 4 2 9 3 10 11 
9 1 5 6 4 3 2 7 8 9 
8 3 2 4 1 5 6 8 7 
14 1 5 3 2 4 6 7 8 9 3 2 3 3 10 
14 1 5 6 7 4 3 2 8 9 2 3 9 3 10 
13 1 5 6 3 2 4 8 7 9 2 3 10 11 
10 1 5 2 3 4 6 7 8 9 10 
14 1 5 6 2 3 4 8 9 7 2 3 3 2 10 
19 1 5 6 7 3 2 4 8 9 2 3 3 2 2 3 10 11 3 2 
13 1 7 5 6 8 4 2 3 9 3 2 10 11 
9 1 5 6 7 2 4 3 8 9 
8 1 5 6 2 4 3 7 8 
30 1 5 6 7 3 4 2 8 9 3 2 3 3 12 2 3 4 2 4 2 3 2 4 2 2 2 2 2 2 13 
21 1 5 6 4 3 2 7 8 9 3 2 9 2 3 2 3 2 3 3 2 10 
51 1 5 6 2 4 3 8 12 3 4 2 2 2 2 2 3 4 2 3 4 4 3 2 9 2 3 2 3 2 3 3 2 2 3 2 3 3 2 2 3 2 3 2 3 2 3 2 3 2 3 10 
20 1 5 3 4 2 6 7 8 9 9 2 3 3 2 3 2 2 3 15 11 
10 1 5 6 4 2 3 7 8 9 10 
7 1 2 3 5 6 7 8 
6 1 5 6 2 3 4 
10 1 5 6 8 3 2 4 9 10 11 
13 1 5 3 2 4 9 6 7 8 9 2 3 10 
3 1 5 6 
8 1 5 6 4 3 2 7 8 
7 1 5 6 3 2 7 8 
12 1 5 6 2 3 4 7 8 9 3 2 10 
10 1 5 6 4 2 3 7 8 9 10 
18 1 5 6 7 8 3 2 4 12 4 3 2 3 2 4 9 10 11 
13 1 5 6 2 3 8 9 3 3 3 3 10 11 
21 2 3 1 5 6 7 8 3 2 4 9 2 4 9 2 3 12 4 2 3 13 
18 1 5 6 4 3 2 8 9 3 2 9 3 2 2 3 2 3 10 
10 1 5 6 2 3 9 9 2 3 10 
6 1 5 6 2 3 4 
3 1 5 6 
10 1 5 6 4 2 3 7 8 9 10 
8 1 5 6 7 4 2 3 8 
8 1 5 6 2 3 4 7 8 
8 1 5 6 2 3 9 10 11 
15 1 5 6 7 2 3 4 8 9 9 3 2 3 10 11 
10 1 5 6 3 4 2 7 8 9 10 
13 1 5 2 3 4 6 7 8 9 2 3 10 11 
8 1 5 6 3 2 4 7 8 
7 1 4 2 3 5 6 8 
20 1 5 6 7 8 2 4 3 12 4 3 4 2 4 3 2 9 2 3 10 
8 1 5 6 3 2 4 9 13 
10 1 7 5 6 8 4 2 3 9 13 
16 1 5 6 7 3 4 2 8 9 5 2 3 3 2 10 11 
6 1 5 2 4 3 6 
8 1 5 4 2 3 6 7 8 
16 1 5 6 2 3 4 8 7 9 9 2 3 2 3 2 10 
13 1 5 6 7 8 2 4 3 9 2 3 10 11 
19 1 5 6 2 3 9 12 2 3 4 3 4 2 2 3 4 9 10 11 
12 1 5 6 7 8 2 4 3 9 2 3 10 
13 1 5 6 2 3 4 7 8 9 2 3 10 11 
15 1 5 6 4 2 3 7 8 9 2 3 9 3 2 10 
12 1 3 4 2 5 6 7 8 9 2 3 10 
10 1 5 6 2 3 7 8 9 9 13 
18 1 5 6 7 8 3 4 2 9 2 3 2 2 3 3 2 9 14 
13 1 5 6 7 2 3 4 8 9 9 3 2 10 
11 1 5 6 3 2 4 8 9 3 2 7 
8 1 5 6 4 2 3 7 8 
16 1 5 2 3 4 6 7 8 9 2 3 4 2 3 3 10 
16 1 5 6 7 2 3 4 8 9 9 3 2 2 3 10 11 
8 1 5 6 2 3 4 9 10 
6 1 5 6 2 3 9 
9 5 1 2 3 4 6 9 7 8 
12 1 5 6 7 8 3 4 2 9 2 3 13 
185 1 5 6 7 3 2 4 8 9 2 9 3 4 2 4 3 2 4 12 3 4 2 3 2 4 4 2 3 3 4 2 3 2 4 2 3 4 4 3 2 4 2 3 4 2 4 3 2 4 3 2 4 4 2 3 2 4 3 3 4 2 3 2 4 3 2 4 2 4 3 3 2 4 3 2 4 4 2 3 2 3 4 2 4 3 3 4 2 2 3 4 2 3 4 2 4 3 9 2 3 2 3 3 2 2 3 2 3 3 2 2 3 3 2 2 3 3 2 3 2 2 3 2 3 2 2 3 9 3 2 2 3 2 3 2 3 3 2 3 2 3 2 2 3 3 2 2 3 3 2 2 3 2 3 3 2 2 2 3 2 3 2 3 3 2 3 2 2 3 2 3 3 2 2 3 2 3 3 2 2 3 2 3 2 14 
13 1 5 6 7 4 2 3 8 9 9 3 2 10 
23 1 5 6 7 8 4 2 3 9 9 12 2 3 4 4 4 2 3 9 2 3 10 11 
7 1 5 6 3 4 2 8 
14 1 5 6 7 3 2 4 8 9 2 3 2 3 10 
16 1 5 3 4 2 6 7 8 12 2 3 4 3 2 4 13 
15 1 5 6 7 8 4 2 3 9 9 2 3 2 3 10 
15 1 5 6 4 3 2 8 9 2 3 9 3 2 3 10 
8 1 5 4 2 3 6 7 8 
36 1 5 6 2 3 4 7 8 9 3 12 3 2 4 4 2 3 2 4 3 3 2 4 4 3 2 9 2 3 9 2 3 3 2 15 11 
15 1 3 2 4 5 6 7 8 9 3 2 2 3 10 11 
14 1 5 6 2 3 4 7 8 9 2 3 9 10 11 
29 1 5 6 2 3 4 7 8 9 3 2 2 3 2 3 2 3 2 3 2 3 2 3 3 2 2 3 10 11 
12 1 5 6 7 4 2 3 8 9 2 3 10 
15 1 5 6 7 4 2 3 8 3 2 9 9 3 2 10 
13 1 5 6 3 4 2 8 7 9 2 3 10 11 
8 1 5 6 3 2 9 3 15 
30 1 5 6 3 4 2 7 8 12 3 2 4 4 2 3 4 2 3 2 3 4 2 3 4 9 3 2 3 2 10 
13 1 5 6 3 4 2 8 9 2 3 3 10 11 
14 1 5 6 2 3 4 2 3 4 7 8 9 3 10 
16 1 5 6 4 3 2 7 8 12 4 2 3 9 2 3 10 
16 1 5 6 2 4 3 7 8 9 3 2 2 3 2 3 10 
7 1 5 6 2 9 2 10 
10 1 7 5 6 8 3 2 4 9 10 
13 1 5 6 7 8 3 2 4 9 3 2 9 10 
13 1 5 6 2 3 4 7 8 9 3 3 10 11 
11 1 5 6 3 2 4 7 8 9 9 10 
13 1 5 3 2 4 6 7 8 9 2 3 3 10 
8 1 5 6 3 2 4 7 8 
14 1 5 6 7 4 2 3 8 9 3 2 2 3 10 
9 1 5 6 2 3 9 3 2 10 
17 1 5 6 7 8 2 4 3 12 2 4 3 9 3 2 2 10 
12 1 3 2 4 5 6 7 8 9 3 2 10 
5 1 5 6 2 3 
5 1 5 6 2 3 
12 1 5 6 8 7 2 3 4 9 2 3 10 
12 1 5 2 3 4 6 7 8 12 2 3 4 
16 1 5 4 3 2 6 7 8 9 2 3 3 2 2 3 10 
26 1 5 6 7 8 12 3 2 4 3 2 4 3 4 2 2 3 4 2 3 4 9 2 3 10 11 
17 1 5 3 2 4 6 7 8 9 2 9 2 2 2 2 10 11 
36 7 1 5 6 4 2 3 8 12 4 3 2 2 3 4 2 4 3 3 2 4 3 4 2 4 2 3 3 2 4 9 3 2 2 10 11 
5 1 5 6 2 3 
5 1 5 6 3 2 
12 1 5 6 2 3 4 7 8 9 3 10 11 
13 1 5 6 2 4 3 9 4 2 3 9 9 14 
7 1 5 6 2 4 3 8 
16 1 5 6 3 2 4 8 7 9 2 3 9 3 2 10 11 
13 1 5 6 2 4 3 7 8 9 2 3 3 10 
9 3 2 1 5 6 2 3 7 8 
13 1 5 6 7 2 3 4 8 9 2 3 3 10 
31 1 5 6 3 4 2 7 8 12 4 2 3 4 2 3 4 9 2 3 2 3 3 2 2 3 2 3 2 3 10 11 
13 1 5 6 2 4 3 8 7 9 3 2 10 11 
13 1 5 6 4 3 2 7 8 9 2 3 10 11 
15 1 5 6 2 4 3 8 7 9 9 2 3 3 2 10 
45 1 5 6 2 3 4 7 8 9 2 3 9 2 3 3 3 2 2 3 2 12 2 3 4 2 2 2 4 2 3 2 2 2 2 3 4 2 2 3 4 9 2 3 10 11 
16 1 5 6 8 7 2 3 4 9 3 2 9 3 2 10 11 
13 1 5 6 2 4 3 7 8 9 9 3 2 10 
8 1 2 3 4 7 5 6 8 
15 1 5 6 2 3 9 9 2 3 3 2 2 2 3 10 
13 1 3 2 4 5 6 7 8 9 3 2 3 10 
36 1 5 6 2 3 4 8 7 12 3 2 4 2 4 4 3 2 2 3 4 2 4 3 4 2 3 9 2 3 2 2 3 2 3 2 10 
5 1 5 2 3 6 
5 1 5 6 3 2 
52 1 5 6 3 2 4 8 7 9 4 3 2 12 2 3 4 9 3 2 2 3 2 3 2 3 2 3 2 3 2 3 2 3 2 3 3 2 2 3 3 2 2 3 3 2 3 2 9 2 3 10 11 
8 1 5 6 3 2 4 7 8 
5 1 3 2 5 6 
17 1 5 6 2 3 4 8 9 7 2 3 3 2 9 9 10 11 
8 1 5 6 2 3 9 3 10 
9 1 5 6 3 2 4 9 10 11 
9 1 3 2 4 5 6 8 9 10 
16 1 5 6 2 3 4 7 8 9 2 3 3 2 2 3 10 
19 1 5 4 2 3 6 7 8 9 4 3 2 9 2 3 3 2 10 11 
13 1 5 6 3 4 2 7 8 9 9 3 2 10 
11 1 5 6 4 2 3 8 7 9 2 3 
9 1 5 6 2 3 4 9 3 10 
5 2 3 1 5 6 
8 1 5 6 4 3 2 7 8 
8 1 5 6 2 3 8 2 3 
16 1 5 6 2 4 3 7 8 9 9 3 2 9 3 2 10 
3 1 5 6 
8 1 5 6 7 8 4 3 2 
9 1 4 2 3 5 6 7 8 2 
8 1 5 6 2 4 3 7 8 
12 1 5 6 8 3 4 2 9 2 3 10 11 
27 1 5 6 7 2 3 4 8 9 3 2 2 3 3 2 2 2 2 2 3 2 3 2 3 2 2 10 
8 1 5 6 7 8 2 4 3 
3 1 5 6 
18 7 1 5 6 3 4 2 8 9 3 3 2 3 2 3 2 3 14 
20 1 5 6 4 2 3 7 8 9 3 2 2 3 2 3 3 2 2 3 10 
12 1 4 2 3 7 5 6 8 9 3 2 10 
23 1 5 6 2 3 4 7 8 9 2 2 3 3 2 3 2 2 3 2 3 2 3 10 
3 1 5 6 
19 1 5 6 2 3 4 4 7 8 9 2 3 9 3 2 3 2 10 11 
17 1 5 6 7 4 2 3 8 9 3 4 2 2 2 3 4 10 
14 1 5 2 4 3 6 7 8 9 9 2 3 10 11 
14 1 5 6 7 3 2 4 8 9 3 2 3 2 10 
11 1 5 6 2 3 4 9 2 3 9 10 
6 1 5 6 3 4 2 
19 1 5 6 3 4 2 7 8 9 2 9 3 3 2 2 2 2 3 15 
8 1 5 7 2 3 4 6 8 
13 1 5 6 7 4 3 2 8 9 2 3 3 13 
14 1 5 6 4 3 2 7 8 12 2 4 3 9 10 
24 1 5 6 2 3 4 7 8 9 2 3 2 3 3 2 2 3 2 3 2 3 10 2 11 
52 1 5 6 3 2 7 8 9 2 3 12 3 4 2 3 4 2 2 3 4 2 4 3 4 3 2 3 2 4 4 2 3 4 3 2 2 3 4 2 3 4 3 2 4 4 2 3 2 4 3 9 10 
10 1 5 7 3 2 4 6 8 9 10 
12 1 5 6 2 3 4 7 8 9 2 3 10 
15 1 5 2 4 3 6 8 9 9 2 3 3 2 10 11 
14 1 5 6 2 3 4 7 8 2 9 3 2 10 11 
10 1 5 6 4 2 3 9 3 2 10 
3 1 5 6 
13 1 5 6 4 3 2 8 9 4 7 2 3 10 
17 1 5 6 3 4 2 7 8 9 9 3 3 2 2 3 9 10 
14 1 5 6 2 3 4 7 8 9 2 9 3 2 15 
18 1 5 6 7 2 3 4 8 9 12 4 2 3 4 3 2 9 13 
13 1 5 6 7 3 2 4 8 9 2 3 10 11 
43 1 5 6 4 2 3 7 8 12 2 4 3 9 2 3 2 3 2 3 2 3 2 2 2 2 2 2 2 2 2 3 2 2 2 2 2 2 2 3 2 2 3 10 
16 1 7 5 6 8 2 4 3 9 2 4 3 2 3 10 11 
11 1 5 6 7 8 3 4 2 9 2 10 
20 1 5 6 4 2 3 7 8 9 2 2 3 2 3 2 3 2 3 10 11 
8 1 5 2 3 4 6 7 8 
8 1 5 4 2 3 6 7 8 
20 1 5 4 2 3 6 7 8 9 9 2 3 9 2 2 3 2 2 3 10 
5 1 5 2 3 6 
14 1 5 6 8 3 2 4 9 9 3 2 3 2 10 
16 1 5 6 4 2 3 7 8 12 2 4 3 9 2 3 10 
12 1 5 6 2 4 3 7 8 9 9 10 11 
25 1 5 2 3 4 6 7 8 9 2 2 3 2 3 2 3 3 2 3 3 2 2 2 3 10 
14 1 5 6 4 2 3 7 8 9 2 2 2 3 10 
5 1 5 6 3 2 
5 1 5 6 2 3 
5 1 5 6 3 2 
12 1 5 6 2 3 4 7 8 9 3 10 11 
25 1 5 6 4 2 3 7 8 9 9 3 2 2 3 2 3 2 3 3 2 3 3 2 10 11 
7 5 1 2 3 4 6 8 
22 1 5 6 3 2 4 8 9 2 3 2 3 3 2 2 3 2 3 3 3 14 11 
24 1 5 6 7 4 2 3 8 9 2 3 2 3 3 2 3 2 2 3 2 3 3 2 10 
8 1 5 6 2 3 4 7 8 
15 1 7 5 2 3 4 6 8 9 3 2 2 3 9 10 
8 1 5 6 7 8 2 3 4 
14 1 5 6 3 2 9 3 2 9 2 3 3 10 11 
8 1 5 6 2 4 3 7 8 
61 1 5 6 3 2 12 3 2 4 2 4 3 4 3 2 2 3 4 3 2 4 2 3 4 2 3 4 2 3 4 4 3 2 9 2 3 4 2 2 3 4 3 2 3 9 3 2 3 2 3 2 2 3 2 3 3 2 2 3 10 11 
11 1 5 6 4 3 2 7 8 9 10 11 
9 1 5 6 2 3 9 2 3 10 
12 1 5 6 2 4 3 7 8 9 3 10 11 
8 1 5 6 3 2 4 8 9 
3 1 5 6 
17 1 5 6 4 3 2 8 7 9 3 2 2 3 2 3 10 11 
13 1 3 4 2 5 6 7 8 9 9 9 10 11 
13 1 5 6 2 3 9 9 3 2 3 2 3 10 
3 1 5 6 
5 1 5 3 2 6 
17 6 1 5 7 8 3 2 4 9 3 2 9 2 3 2 3 10 
20 1 5 6 7 3 2 4 8 9 2 3 3 2 2 3 3 2 2 3 15 
6 1 5 6 2 9 10 
8 1 5 3 2 4 6 7 8 
21 1 5 6 7 8 2 4 3 9 2 3 2 3 9 2 3 2 3 9 9 10 
26 6 1 5 7 8 3 4 2 12 4 2 3 4 2 3 4 2 3 4 9 3 2 3 2 10 11 
14 1 5 6 2 3 4 7 8 9 3 2 2 3 10 
18 1 2 3 4 5 6 7 8 9 3 2 3 9 2 3 3 2 10 
16 1 5 6 3 2 7 8 12 9 2 3 2 3 2 3 10 
10 1 5 6 7 3 2 4 8 9 10 
14 3 2 1 5 6 4 2 3 7 8 9 3 2 10 
3 1 5 6 
5 1 5 6 2 3 
3 1 5 6 
10 1 5 6 2 3 9 2 3 10 11 
66 7 1 5 6 2 4 3 8 4 12 4 3 4 2 4 2 3 2 4 4 3 2 2 4 3 2 3 4 2 3 4 2 3 4 9 2 3 2 3 3 2 3 2 2 3 2 3 2 3 2 3 3 2 2 3 2 2 3 2 3 12 4 2 3 2 13 
9 1 5 6 3 2 9 2 3 10 
7 1 5 6 3 2 9 10 
17 1 5 6 2 3 9 2 2 3 3 2 2 3 2 3 10 11 
8 1 5 6 2 3 4 7 8 
5 1 5 6 3 2 
9 1 5 6 3 4 2 8 9 7 
25 1 5 6 7 3 4 2 8 12 3 2 4 3 4 2 12 2 3 4 2 2 3 4 9 10 
30 1 5 6 2 3 4 8 12 3 2 4 4 2 2 3 4 2 3 4 4 2 3 9 3 2 3 3 2 3 10 
3 1 5 6 
3 1 5 6 
15 1 5 6 2 4 3 7 8 9 3 2 4 2 3 10 
3 1 5 6 
